VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO matrix_multiply
  CLASS BLOCK ;
  FOREIGN matrix_multiply ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 396.000 125.490 400.000 ;
    END
  END clk
  PIN execute
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 396.000 75.810 400.000 ;
    END
  END execute
  PIN input_val[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END input_val[0]
  PIN input_val[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END input_val[1]
  PIN input_val[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END input_val[2]
  PIN input_val[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END input_val[3]
  PIN input_val[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END input_val[4]
  PIN input_val[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END input_val[5]
  PIN input_val[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END input_val[6]
  PIN input_val[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END input_val[7]
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END out[0]
  PIN out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END out[10]
  PIN out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END out[11]
  PIN out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END out[12]
  PIN out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END out[13]
  PIN out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END out[14]
  PIN out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END out[15]
  PIN out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END out[16]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END out[8]
  PIN out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END out[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 396.000 26.130 400.000 ;
    END
  END reset
  PIN sel_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 396.000 175.170 400.000 ;
    END
  END sel_in[0]
  PIN sel_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 396.000 224.850 400.000 ;
    END
  END sel_in[1]
  PIN sel_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 396.000 274.530 400.000 ;
    END
  END sel_in[2]
  PIN sel_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 396.000 324.210 400.000 ;
    END
  END sel_out[0]
  PIN sel_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 396.000 373.890 400.000 ;
    END
  END sel_out[1]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 389.200 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 387.545 394.410 389.150 ;
        RECT 5.330 382.105 394.410 384.935 ;
        RECT 5.330 376.665 394.410 379.495 ;
        RECT 5.330 371.225 394.410 374.055 ;
        RECT 5.330 365.785 394.410 368.615 ;
        RECT 5.330 360.345 394.410 363.175 ;
        RECT 5.330 354.905 394.410 357.735 ;
        RECT 5.330 349.465 394.410 352.295 ;
        RECT 5.330 344.025 394.410 346.855 ;
        RECT 5.330 338.585 394.410 341.415 ;
        RECT 5.330 333.145 394.410 335.975 ;
        RECT 5.330 327.705 394.410 330.535 ;
        RECT 5.330 322.265 394.410 325.095 ;
        RECT 5.330 316.825 394.410 319.655 ;
        RECT 5.330 311.385 394.410 314.215 ;
        RECT 5.330 305.945 394.410 308.775 ;
        RECT 5.330 300.505 394.410 303.335 ;
        RECT 5.330 295.065 394.410 297.895 ;
        RECT 5.330 289.625 394.410 292.455 ;
        RECT 5.330 284.185 394.410 287.015 ;
        RECT 5.330 278.745 394.410 281.575 ;
        RECT 5.330 273.305 394.410 276.135 ;
        RECT 5.330 267.865 394.410 270.695 ;
        RECT 5.330 262.425 394.410 265.255 ;
        RECT 5.330 256.985 394.410 259.815 ;
        RECT 5.330 251.545 394.410 254.375 ;
        RECT 5.330 246.105 394.410 248.935 ;
        RECT 5.330 240.665 394.410 243.495 ;
        RECT 5.330 235.225 394.410 238.055 ;
        RECT 5.330 229.785 394.410 232.615 ;
        RECT 5.330 224.345 394.410 227.175 ;
        RECT 5.330 218.905 394.410 221.735 ;
        RECT 5.330 213.465 394.410 216.295 ;
        RECT 5.330 208.025 394.410 210.855 ;
        RECT 5.330 202.585 394.410 205.415 ;
        RECT 5.330 197.145 394.410 199.975 ;
        RECT 5.330 191.705 394.410 194.535 ;
        RECT 5.330 186.265 394.410 189.095 ;
        RECT 5.330 180.825 394.410 183.655 ;
        RECT 5.330 175.385 394.410 178.215 ;
        RECT 5.330 169.945 394.410 172.775 ;
        RECT 5.330 164.505 394.410 167.335 ;
        RECT 5.330 159.065 394.410 161.895 ;
        RECT 5.330 153.625 394.410 156.455 ;
        RECT 5.330 148.185 394.410 151.015 ;
        RECT 5.330 142.745 394.410 145.575 ;
        RECT 5.330 137.305 394.410 140.135 ;
        RECT 5.330 131.865 394.410 134.695 ;
        RECT 5.330 126.425 394.410 129.255 ;
        RECT 5.330 120.985 394.410 123.815 ;
        RECT 5.330 115.545 394.410 118.375 ;
        RECT 5.330 110.105 394.410 112.935 ;
        RECT 5.330 104.665 394.410 107.495 ;
        RECT 5.330 99.225 394.410 102.055 ;
        RECT 5.330 93.785 394.410 96.615 ;
        RECT 5.330 88.345 394.410 91.175 ;
        RECT 5.330 82.905 394.410 85.735 ;
        RECT 5.330 77.465 394.410 80.295 ;
        RECT 5.330 72.025 394.410 74.855 ;
        RECT 5.330 66.585 394.410 69.415 ;
        RECT 5.330 61.145 394.410 63.975 ;
        RECT 5.330 55.705 394.410 58.535 ;
        RECT 5.330 50.265 394.410 53.095 ;
        RECT 5.330 44.825 394.410 47.655 ;
        RECT 5.330 39.385 394.410 42.215 ;
        RECT 5.330 33.945 394.410 36.775 ;
        RECT 5.330 28.505 394.410 31.335 ;
        RECT 5.330 23.065 394.410 25.895 ;
        RECT 5.330 17.625 394.410 20.455 ;
        RECT 5.330 12.185 394.410 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 394.220 389.045 ;
      LAYER met1 ;
        RECT 5.520 10.240 394.220 389.200 ;
      LAYER met2 ;
        RECT 12.060 395.720 25.570 396.000 ;
        RECT 26.410 395.720 75.250 396.000 ;
        RECT 76.090 395.720 124.930 396.000 ;
        RECT 125.770 395.720 174.610 396.000 ;
        RECT 175.450 395.720 224.290 396.000 ;
        RECT 225.130 395.720 273.970 396.000 ;
        RECT 274.810 395.720 323.650 396.000 ;
        RECT 324.490 395.720 373.330 396.000 ;
        RECT 374.170 395.720 387.680 396.000 ;
        RECT 12.060 4.280 387.680 395.720 ;
        RECT 12.610 4.000 27.410 4.280 ;
        RECT 28.250 4.000 43.050 4.280 ;
        RECT 43.890 4.000 58.690 4.280 ;
        RECT 59.530 4.000 74.330 4.280 ;
        RECT 75.170 4.000 89.970 4.280 ;
        RECT 90.810 4.000 105.610 4.280 ;
        RECT 106.450 4.000 121.250 4.280 ;
        RECT 122.090 4.000 136.890 4.280 ;
        RECT 137.730 4.000 152.530 4.280 ;
        RECT 153.370 4.000 168.170 4.280 ;
        RECT 169.010 4.000 183.810 4.280 ;
        RECT 184.650 4.000 199.450 4.280 ;
        RECT 200.290 4.000 215.090 4.280 ;
        RECT 215.930 4.000 230.730 4.280 ;
        RECT 231.570 4.000 246.370 4.280 ;
        RECT 247.210 4.000 262.010 4.280 ;
        RECT 262.850 4.000 277.650 4.280 ;
        RECT 278.490 4.000 293.290 4.280 ;
        RECT 294.130 4.000 308.930 4.280 ;
        RECT 309.770 4.000 324.570 4.280 ;
        RECT 325.410 4.000 340.210 4.280 ;
        RECT 341.050 4.000 355.850 4.280 ;
        RECT 356.690 4.000 371.490 4.280 ;
        RECT 372.330 4.000 387.130 4.280 ;
      LAYER met3 ;
        RECT 13.865 10.715 385.415 389.125 ;
      LAYER met4 ;
        RECT 66.535 17.175 97.440 387.425 ;
        RECT 99.840 17.175 174.240 387.425 ;
        RECT 176.640 17.175 251.040 387.425 ;
        RECT 253.440 17.175 309.745 387.425 ;
  END
END matrix_multiply
END LIBRARY

