// This is the unpowered netlist.
module matrix_multiply (clk,
    execute,
    reset,
    input_val,
    out,
    sel_in,
    sel_out);
 input clk;
 input execute;
 input reset;
 input [7:0] input_val;
 output [16:0] out;
 input [2:0] sel_in;
 input [1:0] sel_out;

 wire \A[0][0] ;
 wire \A[0][1] ;
 wire \A[0][2] ;
 wire \A[0][3] ;
 wire \A[0][4] ;
 wire \A[0][5] ;
 wire \A[0][6] ;
 wire \A[0][7] ;
 wire \A[1][0] ;
 wire \A[1][1] ;
 wire \A[1][2] ;
 wire \A[1][3] ;
 wire \A[1][4] ;
 wire \A[1][5] ;
 wire \A[1][6] ;
 wire \A[1][7] ;
 wire \A[2][0] ;
 wire \A[2][1] ;
 wire \A[2][2] ;
 wire \A[2][3] ;
 wire \A[2][4] ;
 wire \A[2][5] ;
 wire \A[2][6] ;
 wire \A[2][7] ;
 wire \A[3][0] ;
 wire \A[3][1] ;
 wire \A[3][2] ;
 wire \A[3][3] ;
 wire \A[3][4] ;
 wire \A[3][5] ;
 wire \A[3][6] ;
 wire \A[3][7] ;
 wire \B[0][0] ;
 wire \B[0][1] ;
 wire \B[0][2] ;
 wire \B[0][3] ;
 wire \B[0][4] ;
 wire \B[0][5] ;
 wire \B[0][6] ;
 wire \B[0][7] ;
 wire \B[1][0] ;
 wire \B[1][1] ;
 wire \B[1][2] ;
 wire \B[1][3] ;
 wire \B[1][4] ;
 wire \B[1][5] ;
 wire \B[1][6] ;
 wire \B[1][7] ;
 wire \B[2][0] ;
 wire \B[2][1] ;
 wire \B[2][2] ;
 wire \B[2][3] ;
 wire \B[2][4] ;
 wire \B[2][5] ;
 wire \B[2][6] ;
 wire \B[2][7] ;
 wire \B[3][0] ;
 wire \B[3][1] ;
 wire \B[3][2] ;
 wire \B[3][3] ;
 wire \B[3][4] ;
 wire \B[3][5] ;
 wire \B[3][6] ;
 wire \B[3][7] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;

 sky130_fd_sc_hd__clkbuf_8 _3103_ (.A(\B[3][7] ),
    .X(_0674_));
 sky130_fd_sc_hd__buf_6 _3104_ (.A(_0674_),
    .X(_0685_));
 sky130_fd_sc_hd__clkbuf_8 _3105_ (.A(_0685_),
    .X(_0696_));
 sky130_fd_sc_hd__clkbuf_4 _3106_ (.A(net49),
    .X(_0707_));
 sky130_fd_sc_hd__clkbuf_4 _3107_ (.A(_0707_),
    .X(_0718_));
 sky130_fd_sc_hd__clkbuf_4 _3108_ (.A(\B[1][6] ),
    .X(_0729_));
 sky130_fd_sc_hd__clkbuf_4 _3109_ (.A(_0729_),
    .X(_0740_));
 sky130_fd_sc_hd__buf_2 _3110_ (.A(\A[3][6] ),
    .X(_0751_));
 sky130_fd_sc_hd__clkbuf_4 _3111_ (.A(\A[2][0] ),
    .X(_0762_));
 sky130_fd_sc_hd__buf_2 _3112_ (.A(_0762_),
    .X(_0773_));
 sky130_fd_sc_hd__clkbuf_4 _3113_ (.A(\B[3][0] ),
    .X(_0784_));
 sky130_fd_sc_hd__and4_1 _3114_ (.A(_0740_),
    .B(_0751_),
    .C(_0773_),
    .D(_0784_),
    .X(_0795_));
 sky130_fd_sc_hd__clkbuf_4 _3115_ (.A(\A[3][7] ),
    .X(_0806_));
 sky130_fd_sc_hd__clkbuf_4 _3116_ (.A(\A[2][1] ),
    .X(_0817_));
 sky130_fd_sc_hd__a22o_1 _3117_ (.A1(\B[1][7] ),
    .A2(_0762_),
    .B1(_0817_),
    .B2(\B[1][6] ),
    .X(_0828_));
 sky130_fd_sc_hd__nand4_1 _3118_ (.A(\B[1][6] ),
    .B(\B[1][7] ),
    .C(_0762_),
    .D(_0817_),
    .Y(_0839_));
 sky130_fd_sc_hd__nand4_1 _3119_ (.A(_0806_),
    .B(_0784_),
    .C(_0828_),
    .D(_0839_),
    .Y(_0850_));
 sky130_fd_sc_hd__a22o_1 _3120_ (.A1(_0806_),
    .A2(\B[3][0] ),
    .B1(_0828_),
    .B2(_0839_),
    .X(_0861_));
 sky130_fd_sc_hd__clkbuf_4 _3121_ (.A(net47),
    .X(_0872_));
 sky130_fd_sc_hd__clkbuf_4 _3122_ (.A(_0872_),
    .X(_0883_));
 sky130_fd_sc_hd__nand2_1 _3123_ (.A(\B[1][5] ),
    .B(_0883_),
    .Y(_0894_));
 sky130_fd_sc_hd__buf_2 _3124_ (.A(net57),
    .X(_0905_));
 sky130_fd_sc_hd__clkbuf_4 _3125_ (.A(_0905_),
    .X(_0916_));
 sky130_fd_sc_hd__clkbuf_4 _3126_ (.A(\B[1][3] ),
    .X(_0927_));
 sky130_fd_sc_hd__buf_2 _3127_ (.A(\B[1][4] ),
    .X(_0938_));
 sky130_fd_sc_hd__clkbuf_4 _3128_ (.A(_0938_),
    .X(_0949_));
 sky130_fd_sc_hd__buf_2 _3129_ (.A(net58),
    .X(_0960_));
 sky130_fd_sc_hd__buf_4 _3130_ (.A(_0960_),
    .X(_0971_));
 sky130_fd_sc_hd__a22oi_1 _3131_ (.A1(_0916_),
    .A2(_0927_),
    .B1(_0949_),
    .B2(_0971_),
    .Y(_0982_));
 sky130_fd_sc_hd__buf_2 _3132_ (.A(\A[2][2] ),
    .X(_0993_));
 sky130_fd_sc_hd__clkbuf_4 _3133_ (.A(\A[2][3] ),
    .X(_1004_));
 sky130_fd_sc_hd__buf_2 _3134_ (.A(\B[1][3] ),
    .X(_1015_));
 sky130_fd_sc_hd__clkbuf_4 _3135_ (.A(\B[1][4] ),
    .X(_1026_));
 sky130_fd_sc_hd__and4_1 _3136_ (.A(_0993_),
    .B(_1004_),
    .C(_1015_),
    .D(_1026_),
    .X(_1037_));
 sky130_fd_sc_hd__o21bai_1 _3137_ (.A1(_0894_),
    .A2(_0982_),
    .B1_N(_1037_),
    .Y(_1048_));
 sky130_fd_sc_hd__a21o_1 _3138_ (.A1(_0850_),
    .A2(_0861_),
    .B1(_1048_),
    .X(_1059_));
 sky130_fd_sc_hd__nand3_1 _3139_ (.A(_1048_),
    .B(_0850_),
    .C(_0861_),
    .Y(_1070_));
 sky130_fd_sc_hd__a21bo_1 _3140_ (.A1(_0795_),
    .A2(_1059_),
    .B1_N(_1070_),
    .X(_1081_));
 sky130_fd_sc_hd__buf_2 _3141_ (.A(\B[3][1] ),
    .X(_1092_));
 sky130_fd_sc_hd__buf_4 _3142_ (.A(\B[3][2] ),
    .X(_1103_));
 sky130_fd_sc_hd__buf_2 _3143_ (.A(\A[3][6] ),
    .X(_1114_));
 sky130_fd_sc_hd__a22o_1 _3144_ (.A1(\A[3][7] ),
    .A2(_1092_),
    .B1(_1103_),
    .B2(_1114_),
    .X(_1125_));
 sky130_fd_sc_hd__buf_4 _3145_ (.A(\B[3][1] ),
    .X(_1136_));
 sky130_fd_sc_hd__nand4_1 _3146_ (.A(\A[3][7] ),
    .B(_1114_),
    .C(_1136_),
    .D(_1103_),
    .Y(_1147_));
 sky130_fd_sc_hd__buf_2 _3147_ (.A(\A[3][5] ),
    .X(_1158_));
 sky130_fd_sc_hd__and2_1 _3148_ (.A(_1158_),
    .B(\B[3][3] ),
    .X(_1169_));
 sky130_fd_sc_hd__nand3_1 _3149_ (.A(_1125_),
    .B(_1147_),
    .C(_1169_),
    .Y(_1180_));
 sky130_fd_sc_hd__a21o_1 _3150_ (.A1(_1125_),
    .A2(_1147_),
    .B1(_1169_),
    .X(_1191_));
 sky130_fd_sc_hd__buf_4 _3151_ (.A(\B[3][3] ),
    .X(_1202_));
 sky130_fd_sc_hd__buf_2 _3152_ (.A(net51),
    .X(_1213_));
 sky130_fd_sc_hd__nand2_1 _3153_ (.A(_1202_),
    .B(_1213_),
    .Y(_1224_));
 sky130_fd_sc_hd__clkbuf_4 _3154_ (.A(net42),
    .X(_1235_));
 sky130_fd_sc_hd__a22oi_2 _3155_ (.A1(_1114_),
    .A2(_1235_),
    .B1(_1103_),
    .B2(_1158_),
    .Y(_1246_));
 sky130_fd_sc_hd__buf_2 _3156_ (.A(\B[3][2] ),
    .X(_1257_));
 sky130_fd_sc_hd__and4_1 _3157_ (.A(_1114_),
    .B(_1158_),
    .C(_1092_),
    .D(_1257_),
    .X(_1268_));
 sky130_fd_sc_hd__o21bai_1 _3158_ (.A1(_1224_),
    .A2(_1246_),
    .B1_N(_1268_),
    .Y(_1279_));
 sky130_fd_sc_hd__and3_1 _3159_ (.A(_1180_),
    .B(_1191_),
    .C(_1279_),
    .X(_1290_));
 sky130_fd_sc_hd__a21oi_1 _3160_ (.A1(_1180_),
    .A2(_1191_),
    .B1(_1279_),
    .Y(_1301_));
 sky130_fd_sc_hd__buf_4 _3161_ (.A(\B[3][5] ),
    .X(_1312_));
 sky130_fd_sc_hd__buf_2 _3162_ (.A(\A[3][3] ),
    .X(_1323_));
 sky130_fd_sc_hd__buf_4 _3163_ (.A(\B[3][4] ),
    .X(_1334_));
 sky130_fd_sc_hd__a22oi_1 _3164_ (.A1(_1312_),
    .A2(_1323_),
    .B1(_1213_),
    .B2(_1334_),
    .Y(_1345_));
 sky130_fd_sc_hd__and4_1 _3165_ (.A(\B[3][5] ),
    .B(_1323_),
    .C(_1213_),
    .D(\B[3][4] ),
    .X(_1356_));
 sky130_fd_sc_hd__nor2_1 _3166_ (.A(_1345_),
    .B(_1356_),
    .Y(_1367_));
 sky130_fd_sc_hd__nand2_1 _3167_ (.A(\B[3][6] ),
    .B(_0718_),
    .Y(_1378_));
 sky130_fd_sc_hd__xnor2_1 _3168_ (.A(_1367_),
    .B(_1378_),
    .Y(_1389_));
 sky130_fd_sc_hd__or3b_1 _3169_ (.A(_1290_),
    .B(_1301_),
    .C_N(_1389_),
    .X(_1400_));
 sky130_fd_sc_hd__o21bai_1 _3170_ (.A1(_1290_),
    .A2(_1301_),
    .B1_N(_1389_),
    .Y(_1411_));
 sky130_fd_sc_hd__and3_1 _3171_ (.A(_1081_),
    .B(_1400_),
    .C(_1411_),
    .X(_1422_));
 sky130_fd_sc_hd__or3_1 _3172_ (.A(_1268_),
    .B(_1224_),
    .C(_1246_),
    .X(_1433_));
 sky130_fd_sc_hd__o21ai_1 _3173_ (.A1(_1268_),
    .A2(_1246_),
    .B1(_1224_),
    .Y(_1444_));
 sky130_fd_sc_hd__nand2_1 _3174_ (.A(_1323_),
    .B(\B[3][3] ),
    .Y(_1455_));
 sky130_fd_sc_hd__clkbuf_4 _3175_ (.A(\A[3][4] ),
    .X(_1466_));
 sky130_fd_sc_hd__a22oi_2 _3176_ (.A1(_1158_),
    .A2(_1136_),
    .B1(_1103_),
    .B2(_1466_),
    .Y(_1477_));
 sky130_fd_sc_hd__and4_1 _3177_ (.A(_1158_),
    .B(_1092_),
    .C(\B[3][2] ),
    .D(_1466_),
    .X(_1488_));
 sky130_fd_sc_hd__o21bai_1 _3178_ (.A1(_1455_),
    .A2(_1477_),
    .B1_N(_1488_),
    .Y(_1499_));
 sky130_fd_sc_hd__nand3_1 _3179_ (.A(_1433_),
    .B(_1444_),
    .C(_1499_),
    .Y(_1510_));
 sky130_fd_sc_hd__buf_4 _3180_ (.A(net45),
    .X(_1521_));
 sky130_fd_sc_hd__buf_4 _3181_ (.A(_1323_),
    .X(_1532_));
 sky130_fd_sc_hd__buf_4 _3182_ (.A(\B[3][4] ),
    .X(_1543_));
 sky130_fd_sc_hd__a22oi_1 _3183_ (.A1(_1521_),
    .A2(_0707_),
    .B1(_1532_),
    .B2(_1543_),
    .Y(_1554_));
 sky130_fd_sc_hd__and4_1 _3184_ (.A(_1312_),
    .B(_0707_),
    .C(_1323_),
    .D(_1334_),
    .X(_1565_));
 sky130_fd_sc_hd__nor2_1 _3185_ (.A(_1554_),
    .B(_1565_),
    .Y(_1576_));
 sky130_fd_sc_hd__buf_4 _3186_ (.A(\B[3][6] ),
    .X(_1587_));
 sky130_fd_sc_hd__buf_2 _3187_ (.A(\A[3][1] ),
    .X(_1598_));
 sky130_fd_sc_hd__buf_2 _3188_ (.A(_1598_),
    .X(_1609_));
 sky130_fd_sc_hd__nand2_1 _3189_ (.A(_1587_),
    .B(_1609_),
    .Y(_1620_));
 sky130_fd_sc_hd__xnor2_1 _3190_ (.A(_1576_),
    .B(_1620_),
    .Y(_1630_));
 sky130_fd_sc_hd__a21o_1 _3191_ (.A1(_1433_),
    .A2(_1444_),
    .B1(_1499_),
    .X(_1641_));
 sky130_fd_sc_hd__nand3_1 _3192_ (.A(_1510_),
    .B(_1630_),
    .C(_1641_),
    .Y(_1652_));
 sky130_fd_sc_hd__a21oi_1 _3193_ (.A1(_1400_),
    .A2(_1411_),
    .B1(_1081_),
    .Y(_1663_));
 sky130_fd_sc_hd__a211oi_1 _3194_ (.A1(_1510_),
    .A2(_1652_),
    .B1(_1663_),
    .C1(_1422_),
    .Y(_1674_));
 sky130_fd_sc_hd__o21ba_1 _3195_ (.A1(_1345_),
    .A2(_1378_),
    .B1_N(_1356_),
    .X(_1685_));
 sky130_fd_sc_hd__o21ba_1 _3196_ (.A1(_1422_),
    .A2(_1674_),
    .B1_N(_1685_),
    .X(_1696_));
 sky130_fd_sc_hd__or3b_1 _3197_ (.A(_1422_),
    .B(_1674_),
    .C_N(_1685_),
    .X(_1707_));
 sky130_fd_sc_hd__and2b_1 _3198_ (.A_N(_1696_),
    .B(_1707_),
    .X(_1718_));
 sky130_fd_sc_hd__a31o_1 _3199_ (.A1(_0696_),
    .A2(_0718_),
    .A3(_1718_),
    .B1(_1696_),
    .X(_1729_));
 sky130_fd_sc_hd__buf_2 _3200_ (.A(net55),
    .X(_1740_));
 sky130_fd_sc_hd__a22oi_1 _3201_ (.A1(_1312_),
    .A2(_1213_),
    .B1(_1543_),
    .B2(_1740_),
    .Y(_1751_));
 sky130_fd_sc_hd__and4_1 _3202_ (.A(\B[3][5] ),
    .B(_1740_),
    .C(_1213_),
    .D(_1334_),
    .X(_1762_));
 sky130_fd_sc_hd__nor2_1 _3203_ (.A(_1751_),
    .B(_1762_),
    .Y(_1773_));
 sky130_fd_sc_hd__nand2_1 _3204_ (.A(_1587_),
    .B(_1532_),
    .Y(_1784_));
 sky130_fd_sc_hd__xnor2_1 _3205_ (.A(_1773_),
    .B(_1784_),
    .Y(_1795_));
 sky130_fd_sc_hd__clkbuf_4 _3206_ (.A(_1257_),
    .X(_1806_));
 sky130_fd_sc_hd__nand2_1 _3207_ (.A(_0751_),
    .B(_1806_),
    .Y(_1817_));
 sky130_fd_sc_hd__nand2_1 _3208_ (.A(_0806_),
    .B(_1202_),
    .Y(_1828_));
 sky130_fd_sc_hd__a22o_1 _3209_ (.A1(\A[3][7] ),
    .A2(_1103_),
    .B1(_1202_),
    .B2(_1114_),
    .X(_1839_));
 sky130_fd_sc_hd__o21a_1 _3210_ (.A1(_1817_),
    .A2(_1828_),
    .B1(_1839_),
    .X(_1850_));
 sky130_fd_sc_hd__a21boi_2 _3211_ (.A1(_1125_),
    .A2(_1169_),
    .B1_N(_1147_),
    .Y(_1861_));
 sky130_fd_sc_hd__xnor2_1 _3212_ (.A(_1850_),
    .B(_1861_),
    .Y(_1871_));
 sky130_fd_sc_hd__xnor2_1 _3213_ (.A(_1795_),
    .B(_1871_),
    .Y(_1882_));
 sky130_fd_sc_hd__nand2_1 _3214_ (.A(_0839_),
    .B(_0850_),
    .Y(_1893_));
 sky130_fd_sc_hd__clkbuf_4 _3215_ (.A(\B[1][5] ),
    .X(_1904_));
 sky130_fd_sc_hd__clkbuf_4 _3216_ (.A(net43),
    .X(_1915_));
 sky130_fd_sc_hd__a22o_1 _3217_ (.A1(_0927_),
    .A2(_1915_),
    .B1(_1026_),
    .B2(_1004_),
    .X(_1926_));
 sky130_fd_sc_hd__and4_1 _3218_ (.A(_1004_),
    .B(_1015_),
    .C(_1915_),
    .D(_0938_),
    .X(_1937_));
 sky130_fd_sc_hd__a31oi_2 _3219_ (.A1(_1904_),
    .A2(_0971_),
    .A3(_1926_),
    .B1(_1937_),
    .Y(_1948_));
 sky130_fd_sc_hd__clkbuf_4 _3220_ (.A(\B[1][7] ),
    .X(_1959_));
 sky130_fd_sc_hd__a22oi_2 _3221_ (.A1(_1959_),
    .A2(_0883_),
    .B1(_0971_),
    .B2(_0729_),
    .Y(_1970_));
 sky130_fd_sc_hd__and4_1 _3222_ (.A(_0729_),
    .B(\B[1][7] ),
    .C(_0817_),
    .D(_0971_),
    .X(_1981_));
 sky130_fd_sc_hd__nor2_1 _3223_ (.A(_1970_),
    .B(_1981_),
    .Y(_1992_));
 sky130_fd_sc_hd__xnor2_1 _3224_ (.A(_1948_),
    .B(_1992_),
    .Y(_2003_));
 sky130_fd_sc_hd__or3_1 _3225_ (.A(_1948_),
    .B(_1970_),
    .C(_1981_),
    .X(_2014_));
 sky130_fd_sc_hd__a21bo_1 _3226_ (.A1(_1893_),
    .A2(_2003_),
    .B1_N(_2014_),
    .X(_2024_));
 sky130_fd_sc_hd__and2b_1 _3227_ (.A_N(_1882_),
    .B(_2024_),
    .X(_2035_));
 sky130_fd_sc_hd__nor3b_1 _3228_ (.A(_1290_),
    .B(_1301_),
    .C_N(_1389_),
    .Y(_2046_));
 sky130_fd_sc_hd__xnor2_1 _3229_ (.A(_2024_),
    .B(_1882_),
    .Y(_2057_));
 sky130_fd_sc_hd__o21a_1 _3230_ (.A1(_1290_),
    .A2(_2046_),
    .B1(_2057_),
    .X(_2068_));
 sky130_fd_sc_hd__o21ba_1 _3231_ (.A1(_1751_),
    .A2(_1784_),
    .B1_N(_1762_),
    .X(_2079_));
 sky130_fd_sc_hd__o21ba_1 _3232_ (.A1(_2035_),
    .A2(_2068_),
    .B1_N(_2079_),
    .X(_2090_));
 sky130_fd_sc_hd__or3b_1 _3233_ (.A(_2035_),
    .B(_2068_),
    .C_N(_2079_),
    .X(_2101_));
 sky130_fd_sc_hd__and2b_1 _3234_ (.A_N(_2090_),
    .B(_2101_),
    .X(_2112_));
 sky130_fd_sc_hd__nand2_1 _3235_ (.A(\B[3][7] ),
    .B(_1532_),
    .Y(_2123_));
 sky130_fd_sc_hd__xnor2_1 _3236_ (.A(_2112_),
    .B(_2123_),
    .Y(_2133_));
 sky130_fd_sc_hd__inv_2 _3237_ (.A(_1839_),
    .Y(_2144_));
 sky130_fd_sc_hd__nor2_2 _3238_ (.A(_1817_),
    .B(_1828_),
    .Y(_2155_));
 sky130_fd_sc_hd__nand2_1 _3239_ (.A(_1795_),
    .B(_1871_),
    .Y(_2166_));
 sky130_fd_sc_hd__o31ai_4 _3240_ (.A1(_2144_),
    .A2(_2155_),
    .A3(_1861_),
    .B1(_2166_),
    .Y(_2177_));
 sky130_fd_sc_hd__a22oi_1 _3241_ (.A1(\B[1][7] ),
    .A2(_0971_),
    .B1(_0916_),
    .B2(_0729_),
    .Y(_2188_));
 sky130_fd_sc_hd__and4_1 _3242_ (.A(\B[1][6] ),
    .B(\B[1][7] ),
    .C(_0993_),
    .D(_1004_),
    .X(_2198_));
 sky130_fd_sc_hd__or2_1 _3243_ (.A(_2188_),
    .B(_2198_),
    .X(_2208_));
 sky130_fd_sc_hd__clkbuf_4 _3244_ (.A(net50),
    .X(_2218_));
 sky130_fd_sc_hd__a22o_1 _3245_ (.A1(_2218_),
    .A2(_1015_),
    .B1(_1915_),
    .B2(_0938_),
    .X(_2228_));
 sky130_fd_sc_hd__clkbuf_4 _3246_ (.A(\A[2][4] ),
    .X(_2238_));
 sky130_fd_sc_hd__and4_1 _3247_ (.A(_2218_),
    .B(_1015_),
    .C(_2238_),
    .D(_0938_),
    .X(_2248_));
 sky130_fd_sc_hd__a31o_1 _3248_ (.A1(_1904_),
    .A2(_0916_),
    .A3(_2228_),
    .B1(_2248_),
    .X(_2259_));
 sky130_fd_sc_hd__or2b_1 _3249_ (.A(_2208_),
    .B_N(_2259_),
    .X(_2269_));
 sky130_fd_sc_hd__xnor2_1 _3250_ (.A(_2259_),
    .B(_2208_),
    .Y(_2279_));
 sky130_fd_sc_hd__nand2_1 _3251_ (.A(_1981_),
    .B(_2279_),
    .Y(_2289_));
 sky130_fd_sc_hd__and3_1 _3252_ (.A(\B[3][5] ),
    .B(_0751_),
    .C(_1740_),
    .X(_2300_));
 sky130_fd_sc_hd__a22o_1 _3253_ (.A1(\B[3][5] ),
    .A2(_1740_),
    .B1(_1334_),
    .B2(_0751_),
    .X(_2310_));
 sky130_fd_sc_hd__a21bo_1 _3254_ (.A1(_1543_),
    .A2(_2300_),
    .B1_N(_2310_),
    .X(_2320_));
 sky130_fd_sc_hd__nand2_1 _3255_ (.A(_1587_),
    .B(_1213_),
    .Y(_2330_));
 sky130_fd_sc_hd__xor2_1 _3256_ (.A(_2320_),
    .B(_2330_),
    .X(_2340_));
 sky130_fd_sc_hd__clkbuf_4 _3257_ (.A(_1202_),
    .X(_2347_));
 sky130_fd_sc_hd__and3_1 _3258_ (.A(_0806_),
    .B(_2347_),
    .C(_1817_),
    .X(_2354_));
 sky130_fd_sc_hd__xnor2_1 _3259_ (.A(_2340_),
    .B(_2354_),
    .Y(_2360_));
 sky130_fd_sc_hd__a21oi_1 _3260_ (.A1(_2269_),
    .A2(_2289_),
    .B1(_2360_),
    .Y(_2367_));
 sky130_fd_sc_hd__nand3_1 _3261_ (.A(_2269_),
    .B(_2289_),
    .C(_2360_),
    .Y(_2373_));
 sky130_fd_sc_hd__and2b_1 _3262_ (.A_N(_2367_),
    .B(_2373_),
    .X(_2379_));
 sky130_fd_sc_hd__xor2_2 _3263_ (.A(_2177_),
    .B(_2379_),
    .X(_2385_));
 sky130_fd_sc_hd__clkbuf_4 _3264_ (.A(\A[2][6] ),
    .X(_2392_));
 sky130_fd_sc_hd__a22o_1 _3265_ (.A1(_2392_),
    .A2(_1015_),
    .B1(_0938_),
    .B2(_2218_),
    .X(_2399_));
 sky130_fd_sc_hd__clkbuf_4 _3266_ (.A(\A[2][6] ),
    .X(_2405_));
 sky130_fd_sc_hd__nand4_1 _3267_ (.A(_2405_),
    .B(_2218_),
    .C(_0927_),
    .D(_1026_),
    .Y(_2411_));
 sky130_fd_sc_hd__and2_1 _3268_ (.A(\B[1][5] ),
    .B(_2238_),
    .X(_2417_));
 sky130_fd_sc_hd__a21o_1 _3269_ (.A1(_2399_),
    .A2(_2411_),
    .B1(_2417_),
    .X(_2424_));
 sky130_fd_sc_hd__nand3_1 _3270_ (.A(_2399_),
    .B(_2411_),
    .C(_2417_),
    .Y(_2430_));
 sky130_fd_sc_hd__clkbuf_4 _3271_ (.A(\A[2][7] ),
    .X(_2431_));
 sky130_fd_sc_hd__clkbuf_4 _3272_ (.A(net41),
    .X(_2432_));
 sky130_fd_sc_hd__buf_4 _3273_ (.A(net44),
    .X(_2433_));
 sky130_fd_sc_hd__nand2_1 _3274_ (.A(_2405_),
    .B(_2433_),
    .Y(_2434_));
 sky130_fd_sc_hd__and3_1 _3275_ (.A(_2431_),
    .B(_2432_),
    .C(_2434_),
    .X(_2435_));
 sky130_fd_sc_hd__and3_2 _3276_ (.A(_2424_),
    .B(_2430_),
    .C(_2435_),
    .X(_2436_));
 sky130_fd_sc_hd__clkbuf_4 _3277_ (.A(\B[1][1] ),
    .X(_2437_));
 sky130_fd_sc_hd__clkbuf_4 _3278_ (.A(\B[1][2] ),
    .X(_2438_));
 sky130_fd_sc_hd__and4_1 _3279_ (.A(\A[2][7] ),
    .B(_2392_),
    .C(_2437_),
    .D(_2438_),
    .X(_2439_));
 sky130_fd_sc_hd__clkbuf_4 _3280_ (.A(_1015_),
    .X(_2440_));
 sky130_fd_sc_hd__nand2_1 _3281_ (.A(_2431_),
    .B(_2440_),
    .Y(_2441_));
 sky130_fd_sc_hd__nand2_1 _3282_ (.A(_2405_),
    .B(_1026_),
    .Y(_2442_));
 sky130_fd_sc_hd__and4_1 _3283_ (.A(_2431_),
    .B(_2405_),
    .C(_0927_),
    .D(_1026_),
    .X(_2443_));
 sky130_fd_sc_hd__a21oi_1 _3284_ (.A1(_2441_),
    .A2(_2442_),
    .B1(_2443_),
    .Y(_2444_));
 sky130_fd_sc_hd__clkbuf_4 _3285_ (.A(_2218_),
    .X(_2445_));
 sky130_fd_sc_hd__nand2_1 _3286_ (.A(_1904_),
    .B(_2445_),
    .Y(_2446_));
 sky130_fd_sc_hd__xnor2_1 _3287_ (.A(_2444_),
    .B(_2446_),
    .Y(_2447_));
 sky130_fd_sc_hd__o21a_1 _3288_ (.A1(_2436_),
    .A2(_2439_),
    .B1(_2447_),
    .X(_2448_));
 sky130_fd_sc_hd__or3_1 _3289_ (.A(_2447_),
    .B(_2436_),
    .C(_2439_),
    .X(_2449_));
 sky130_fd_sc_hd__and2b_1 _3290_ (.A_N(_2448_),
    .B(_2449_),
    .X(_2450_));
 sky130_fd_sc_hd__a21bo_1 _3291_ (.A1(_2399_),
    .A2(_2417_),
    .B1_N(_2411_),
    .X(_2451_));
 sky130_fd_sc_hd__nand2_1 _3292_ (.A(_1959_),
    .B(_0916_),
    .Y(_2452_));
 sky130_fd_sc_hd__nand2_1 _3293_ (.A(_0729_),
    .B(_1915_),
    .Y(_2453_));
 sky130_fd_sc_hd__and4_1 _3294_ (.A(_0729_),
    .B(\B[1][7] ),
    .C(_1004_),
    .D(_1915_),
    .X(_2454_));
 sky130_fd_sc_hd__a21o_1 _3295_ (.A1(_2452_),
    .A2(_2453_),
    .B1(_2454_),
    .X(_2455_));
 sky130_fd_sc_hd__xnor2_1 _3296_ (.A(_2451_),
    .B(_2455_),
    .Y(_2456_));
 sky130_fd_sc_hd__nor2_1 _3297_ (.A(_2198_),
    .B(_2456_),
    .Y(_2457_));
 sky130_fd_sc_hd__and2_1 _3298_ (.A(_2198_),
    .B(_2456_),
    .X(_2458_));
 sky130_fd_sc_hd__nor2_1 _3299_ (.A(_2457_),
    .B(_2458_),
    .Y(_2459_));
 sky130_fd_sc_hd__xor2_2 _3300_ (.A(_2450_),
    .B(_2459_),
    .X(_2460_));
 sky130_fd_sc_hd__a21oi_2 _3301_ (.A1(_2424_),
    .A2(_2430_),
    .B1(_2435_),
    .Y(_2461_));
 sky130_fd_sc_hd__and2b_1 _3302_ (.A_N(_2248_),
    .B(_2228_),
    .X(_2462_));
 sky130_fd_sc_hd__nand2_1 _3303_ (.A(_1904_),
    .B(_0916_),
    .Y(_2463_));
 sky130_fd_sc_hd__xnor2_1 _3304_ (.A(_2462_),
    .B(_2463_),
    .Y(_2464_));
 sky130_fd_sc_hd__a22oi_1 _3305_ (.A1(_2431_),
    .A2(_2433_),
    .B1(_2432_),
    .B2(_2405_),
    .Y(_2465_));
 sky130_fd_sc_hd__or2_1 _3306_ (.A(_2439_),
    .B(_2465_),
    .X(_2466_));
 sky130_fd_sc_hd__and2_1 _3307_ (.A(_2218_),
    .B(_2438_),
    .X(_2467_));
 sky130_fd_sc_hd__clkbuf_4 _3308_ (.A(\B[1][0] ),
    .X(_2468_));
 sky130_fd_sc_hd__a22o_1 _3309_ (.A1(\A[2][7] ),
    .A2(_2468_),
    .B1(_2437_),
    .B2(_2405_),
    .X(_2469_));
 sky130_fd_sc_hd__clkbuf_4 _3310_ (.A(\B[1][0] ),
    .X(_2470_));
 sky130_fd_sc_hd__buf_4 _3311_ (.A(_2470_),
    .X(_2471_));
 sky130_fd_sc_hd__nand4_2 _3312_ (.A(_2431_),
    .B(_2405_),
    .C(_2471_),
    .D(_2433_),
    .Y(_2472_));
 sky130_fd_sc_hd__a21bo_1 _3313_ (.A1(_2467_),
    .A2(_2469_),
    .B1_N(_2472_),
    .X(_2473_));
 sky130_fd_sc_hd__xnor2_1 _3314_ (.A(_2466_),
    .B(_2473_),
    .Y(_2474_));
 sky130_fd_sc_hd__or2b_1 _3315_ (.A(_2466_),
    .B_N(_2473_),
    .X(_2475_));
 sky130_fd_sc_hd__a21boi_2 _3316_ (.A1(_2464_),
    .A2(_2474_),
    .B1_N(_2475_),
    .Y(_2476_));
 sky130_fd_sc_hd__or2_1 _3317_ (.A(_1981_),
    .B(_2279_),
    .X(_2477_));
 sky130_fd_sc_hd__nand2_2 _3318_ (.A(_2289_),
    .B(_2477_),
    .Y(_2478_));
 sky130_fd_sc_hd__or2_1 _3319_ (.A(_2436_),
    .B(_2461_),
    .X(_2479_));
 sky130_fd_sc_hd__xnor2_2 _3320_ (.A(_2479_),
    .B(_2476_),
    .Y(_2480_));
 sky130_fd_sc_hd__o32ai_4 _3321_ (.A1(_2436_),
    .A2(_2461_),
    .A3(_2476_),
    .B1(_2478_),
    .B2(_2480_),
    .Y(_2481_));
 sky130_fd_sc_hd__xor2_2 _3322_ (.A(_2460_),
    .B(_2481_),
    .X(_2482_));
 sky130_fd_sc_hd__xnor2_2 _3323_ (.A(_2385_),
    .B(_2482_),
    .Y(_2483_));
 sky130_fd_sc_hd__nor3_1 _3324_ (.A(_1290_),
    .B(_2046_),
    .C(_2057_),
    .Y(_2484_));
 sky130_fd_sc_hd__nor2_1 _3325_ (.A(_2068_),
    .B(_2484_),
    .Y(_2485_));
 sky130_fd_sc_hd__xor2_2 _3326_ (.A(_2478_),
    .B(_2480_),
    .X(_2486_));
 sky130_fd_sc_hd__xnor2_2 _3327_ (.A(_1893_),
    .B(_2003_),
    .Y(_2487_));
 sky130_fd_sc_hd__xnor2_1 _3328_ (.A(_2464_),
    .B(_2474_),
    .Y(_2488_));
 sky130_fd_sc_hd__nand2_1 _3329_ (.A(_1904_),
    .B(_0971_),
    .Y(_2489_));
 sky130_fd_sc_hd__and2b_1 _3330_ (.A_N(_1937_),
    .B(_1926_),
    .X(_2490_));
 sky130_fd_sc_hd__xnor2_1 _3331_ (.A(_2489_),
    .B(_2490_),
    .Y(_2491_));
 sky130_fd_sc_hd__nand3_1 _3332_ (.A(_2472_),
    .B(_2467_),
    .C(_2469_),
    .Y(_2492_));
 sky130_fd_sc_hd__a21o_1 _3333_ (.A1(_2472_),
    .A2(_2469_),
    .B1(_2467_),
    .X(_2493_));
 sky130_fd_sc_hd__nand2_1 _3334_ (.A(_2438_),
    .B(_1915_),
    .Y(_2494_));
 sky130_fd_sc_hd__a22oi_2 _3335_ (.A1(_2405_),
    .A2(_2468_),
    .B1(_2437_),
    .B2(_2218_),
    .Y(_2495_));
 sky130_fd_sc_hd__clkbuf_4 _3336_ (.A(\B[1][1] ),
    .X(_2496_));
 sky130_fd_sc_hd__and4_1 _3337_ (.A(_2392_),
    .B(_2218_),
    .C(_2470_),
    .D(_2496_),
    .X(_2497_));
 sky130_fd_sc_hd__o21bai_1 _3338_ (.A1(_2494_),
    .A2(_2495_),
    .B1_N(_2497_),
    .Y(_2498_));
 sky130_fd_sc_hd__a21o_1 _3339_ (.A1(_2492_),
    .A2(_2493_),
    .B1(_2498_),
    .X(_2499_));
 sky130_fd_sc_hd__nand3_1 _3340_ (.A(_2492_),
    .B(_2493_),
    .C(_2498_),
    .Y(_2500_));
 sky130_fd_sc_hd__a21bo_1 _3341_ (.A1(_2491_),
    .A2(_2499_),
    .B1_N(_2500_),
    .X(_2501_));
 sky130_fd_sc_hd__xor2_2 _3342_ (.A(_2488_),
    .B(_2501_),
    .X(_2502_));
 sky130_fd_sc_hd__or2b_1 _3343_ (.A(_2488_),
    .B_N(_2501_),
    .X(_2503_));
 sky130_fd_sc_hd__o21a_1 _3344_ (.A1(_2487_),
    .A2(_2502_),
    .B1(_2503_),
    .X(_2504_));
 sky130_fd_sc_hd__xnor2_2 _3345_ (.A(_2486_),
    .B(_2504_),
    .Y(_2505_));
 sky130_fd_sc_hd__or2b_1 _3346_ (.A(_2504_),
    .B_N(_2486_),
    .X(_2506_));
 sky130_fd_sc_hd__a21boi_2 _3347_ (.A1(_2485_),
    .A2(_2505_),
    .B1_N(_2506_),
    .Y(_2507_));
 sky130_fd_sc_hd__xor2_2 _3348_ (.A(_2483_),
    .B(_2507_),
    .X(_2508_));
 sky130_fd_sc_hd__xnor2_2 _3349_ (.A(_2133_),
    .B(_2508_),
    .Y(_2509_));
 sky130_fd_sc_hd__nand2_1 _3350_ (.A(\B[3][7] ),
    .B(_0718_),
    .Y(_2510_));
 sky130_fd_sc_hd__xnor2_1 _3351_ (.A(_1718_),
    .B(_2510_),
    .Y(_2511_));
 sky130_fd_sc_hd__xnor2_1 _3352_ (.A(_2485_),
    .B(_2505_),
    .Y(_2512_));
 sky130_fd_sc_hd__o211a_1 _3353_ (.A1(_1422_),
    .A2(_1663_),
    .B1(_1652_),
    .C1(_1510_),
    .X(_2513_));
 sky130_fd_sc_hd__nor2_1 _3354_ (.A(_1674_),
    .B(_2513_),
    .Y(_2514_));
 sky130_fd_sc_hd__xnor2_2 _3355_ (.A(_2487_),
    .B(_2502_),
    .Y(_2515_));
 sky130_fd_sc_hd__and3_1 _3356_ (.A(_1070_),
    .B(_0795_),
    .C(_1059_),
    .X(_2516_));
 sky130_fd_sc_hd__a21oi_1 _3357_ (.A1(_1070_),
    .A2(_1059_),
    .B1(_0795_),
    .Y(_2517_));
 sky130_fd_sc_hd__or2_1 _3358_ (.A(_2516_),
    .B(_2517_),
    .X(_2518_));
 sky130_fd_sc_hd__nand3_1 _3359_ (.A(_2500_),
    .B(_2491_),
    .C(_2499_),
    .Y(_2519_));
 sky130_fd_sc_hd__a21o_1 _3360_ (.A1(_2500_),
    .A2(_2499_),
    .B1(_2491_),
    .X(_2520_));
 sky130_fd_sc_hd__nor2_1 _3361_ (.A(_1037_),
    .B(_0982_),
    .Y(_2521_));
 sky130_fd_sc_hd__xnor2_1 _3362_ (.A(_0894_),
    .B(_2521_),
    .Y(_2522_));
 sky130_fd_sc_hd__or3_1 _3363_ (.A(_2497_),
    .B(_2494_),
    .C(_2495_),
    .X(_2523_));
 sky130_fd_sc_hd__o21ai_1 _3364_ (.A1(_2497_),
    .A2(_2495_),
    .B1(_2494_),
    .Y(_2524_));
 sky130_fd_sc_hd__nand2_1 _3365_ (.A(_2438_),
    .B(_0905_),
    .Y(_2525_));
 sky130_fd_sc_hd__buf_2 _3366_ (.A(\A[2][5] ),
    .X(_2526_));
 sky130_fd_sc_hd__a22oi_2 _3367_ (.A1(_2526_),
    .A2(_2470_),
    .B1(_2496_),
    .B2(_2238_),
    .Y(_2527_));
 sky130_fd_sc_hd__and4_1 _3368_ (.A(\A[2][5] ),
    .B(\B[1][0] ),
    .C(\B[1][1] ),
    .D(\A[2][4] ),
    .X(_2528_));
 sky130_fd_sc_hd__o21bai_1 _3369_ (.A1(_2525_),
    .A2(_2527_),
    .B1_N(_2528_),
    .Y(_2529_));
 sky130_fd_sc_hd__a21o_1 _3370_ (.A1(_2523_),
    .A2(_2524_),
    .B1(_2529_),
    .X(_2530_));
 sky130_fd_sc_hd__nand3_1 _3371_ (.A(_2523_),
    .B(_2524_),
    .C(_2529_),
    .Y(_2531_));
 sky130_fd_sc_hd__a21bo_1 _3372_ (.A1(_2522_),
    .A2(_2530_),
    .B1_N(_2531_),
    .X(_2532_));
 sky130_fd_sc_hd__a21oi_1 _3373_ (.A1(_2519_),
    .A2(_2520_),
    .B1(_2532_),
    .Y(_2533_));
 sky130_fd_sc_hd__and3_1 _3374_ (.A(_2519_),
    .B(_2520_),
    .C(_2532_),
    .X(_2534_));
 sky130_fd_sc_hd__o21ba_1 _3375_ (.A1(_2518_),
    .A2(_2533_),
    .B1_N(_2534_),
    .X(_2535_));
 sky130_fd_sc_hd__xor2_2 _3376_ (.A(_2515_),
    .B(_2535_),
    .X(_2536_));
 sky130_fd_sc_hd__nor2_1 _3377_ (.A(_2515_),
    .B(_2535_),
    .Y(_2537_));
 sky130_fd_sc_hd__a21o_1 _3378_ (.A1(_2514_),
    .A2(_2536_),
    .B1(_2537_),
    .X(_2538_));
 sky130_fd_sc_hd__xnor2_1 _3379_ (.A(_2512_),
    .B(_2538_),
    .Y(_2539_));
 sky130_fd_sc_hd__or2b_1 _3380_ (.A(_2512_),
    .B_N(_2538_),
    .X(_2540_));
 sky130_fd_sc_hd__a21boi_2 _3381_ (.A1(_2511_),
    .A2(_2539_),
    .B1_N(_2540_),
    .Y(_2541_));
 sky130_fd_sc_hd__xor2_2 _3382_ (.A(_2509_),
    .B(_2541_),
    .X(_2542_));
 sky130_fd_sc_hd__xnor2_2 _3383_ (.A(_1729_),
    .B(_2542_),
    .Y(_2543_));
 sky130_fd_sc_hd__clkbuf_4 _3384_ (.A(_1609_),
    .X(_2544_));
 sky130_fd_sc_hd__and4_1 _3385_ (.A(_0872_),
    .B(\A[2][2] ),
    .C(\B[1][3] ),
    .D(\B[1][4] ),
    .X(_2545_));
 sky130_fd_sc_hd__nand2_1 _3386_ (.A(\B[1][5] ),
    .B(_0762_),
    .Y(_2546_));
 sky130_fd_sc_hd__a22oi_1 _3387_ (.A1(_0993_),
    .A2(_1015_),
    .B1(_0938_),
    .B2(_0872_),
    .Y(_2547_));
 sky130_fd_sc_hd__or2_1 _3388_ (.A(_2547_),
    .B(_2545_),
    .X(_2548_));
 sky130_fd_sc_hd__nor2_1 _3389_ (.A(_2546_),
    .B(_2548_),
    .Y(_2549_));
 sky130_fd_sc_hd__clkbuf_4 _3390_ (.A(_0773_),
    .X(_2550_));
 sky130_fd_sc_hd__buf_2 _3391_ (.A(_0751_),
    .X(_2551_));
 sky130_fd_sc_hd__a22oi_1 _3392_ (.A1(_0740_),
    .A2(_2550_),
    .B1(_0784_),
    .B2(_2551_),
    .Y(_2552_));
 sky130_fd_sc_hd__nor2_1 _3393_ (.A(_0795_),
    .B(_2552_),
    .Y(_2553_));
 sky130_fd_sc_hd__o21a_2 _3394_ (.A1(_2545_),
    .A2(_2549_),
    .B1(_2553_),
    .X(_2554_));
 sky130_fd_sc_hd__a21o_1 _3395_ (.A1(_1510_),
    .A2(_1641_),
    .B1(_1630_),
    .X(_2555_));
 sky130_fd_sc_hd__and3_1 _3396_ (.A(_1652_),
    .B(_2554_),
    .C(_2555_),
    .X(_2556_));
 sky130_fd_sc_hd__or3_1 _3397_ (.A(_1488_),
    .B(_1455_),
    .C(_1477_),
    .X(_2557_));
 sky130_fd_sc_hd__o21ai_1 _3398_ (.A1(_1488_),
    .A2(_1477_),
    .B1(_1455_),
    .Y(_2558_));
 sky130_fd_sc_hd__buf_2 _3399_ (.A(\A[3][2] ),
    .X(_2559_));
 sky130_fd_sc_hd__nand2_1 _3400_ (.A(_2559_),
    .B(\B[3][3] ),
    .Y(_2560_));
 sky130_fd_sc_hd__a22oi_2 _3401_ (.A1(_1257_),
    .A2(\A[3][3] ),
    .B1(_1466_),
    .B2(_1136_),
    .Y(_2561_));
 sky130_fd_sc_hd__and4_1 _3402_ (.A(\B[3][1] ),
    .B(\B[3][2] ),
    .C(\A[3][3] ),
    .D(_1466_),
    .X(_2562_));
 sky130_fd_sc_hd__o21bai_1 _3403_ (.A1(_2560_),
    .A2(_2561_),
    .B1_N(_2562_),
    .Y(_2563_));
 sky130_fd_sc_hd__nand3_1 _3404_ (.A(_2557_),
    .B(_2558_),
    .C(_2563_),
    .Y(_2564_));
 sky130_fd_sc_hd__a22oi_1 _3405_ (.A1(_1312_),
    .A2(_1598_),
    .B1(_0707_),
    .B2(_1334_),
    .Y(_2565_));
 sky130_fd_sc_hd__and4_1 _3406_ (.A(\B[3][5] ),
    .B(_1598_),
    .C(_0707_),
    .D(\B[3][4] ),
    .X(_2566_));
 sky130_fd_sc_hd__nor2_1 _3407_ (.A(_2565_),
    .B(_2566_),
    .Y(_2567_));
 sky130_fd_sc_hd__buf_2 _3408_ (.A(\A[3][0] ),
    .X(_2568_));
 sky130_fd_sc_hd__nand2_1 _3409_ (.A(_1587_),
    .B(_2568_),
    .Y(_2569_));
 sky130_fd_sc_hd__xnor2_1 _3410_ (.A(_2567_),
    .B(_2569_),
    .Y(_2570_));
 sky130_fd_sc_hd__a21o_1 _3411_ (.A1(_2557_),
    .A2(_2558_),
    .B1(_2563_),
    .X(_2571_));
 sky130_fd_sc_hd__nand3_1 _3412_ (.A(_2564_),
    .B(_2570_),
    .C(_2571_),
    .Y(_2572_));
 sky130_fd_sc_hd__nand2_1 _3413_ (.A(_2564_),
    .B(_2572_),
    .Y(_2573_));
 sky130_fd_sc_hd__nand3_1 _3414_ (.A(_1652_),
    .B(_2554_),
    .C(_2555_),
    .Y(_2574_));
 sky130_fd_sc_hd__a21o_1 _3415_ (.A1(_1652_),
    .A2(_2555_),
    .B1(_2554_),
    .X(_2575_));
 sky130_fd_sc_hd__and3_1 _3416_ (.A(_2573_),
    .B(_2574_),
    .C(_2575_),
    .X(_2576_));
 sky130_fd_sc_hd__o21ba_1 _3417_ (.A1(_1554_),
    .A2(_1620_),
    .B1_N(_1565_),
    .X(_2577_));
 sky130_fd_sc_hd__o21ba_1 _3418_ (.A1(_2556_),
    .A2(_2576_),
    .B1_N(_2577_),
    .X(_2578_));
 sky130_fd_sc_hd__or3b_1 _3419_ (.A(_2556_),
    .B(_2576_),
    .C_N(_2577_),
    .X(_2579_));
 sky130_fd_sc_hd__and2b_1 _3420_ (.A_N(_2578_),
    .B(_2579_),
    .X(_2580_));
 sky130_fd_sc_hd__a31o_1 _3421_ (.A1(_0685_),
    .A2(_2544_),
    .A3(_2580_),
    .B1(_2578_),
    .X(_2581_));
 sky130_fd_sc_hd__xor2_1 _3422_ (.A(_2511_),
    .B(_2539_),
    .X(_2582_));
 sky130_fd_sc_hd__nand2_1 _3423_ (.A(_0674_),
    .B(_2544_),
    .Y(_2583_));
 sky130_fd_sc_hd__xor2_2 _3424_ (.A(_2580_),
    .B(_2583_),
    .X(_2584_));
 sky130_fd_sc_hd__xnor2_1 _3425_ (.A(_2514_),
    .B(_2536_),
    .Y(_2585_));
 sky130_fd_sc_hd__a21oi_1 _3426_ (.A1(_2574_),
    .A2(_2575_),
    .B1(_2573_),
    .Y(_2586_));
 sky130_fd_sc_hd__nor2_1 _3427_ (.A(_2576_),
    .B(_2586_),
    .Y(_2587_));
 sky130_fd_sc_hd__or3_1 _3428_ (.A(_2534_),
    .B(_2518_),
    .C(_2533_),
    .X(_2588_));
 sky130_fd_sc_hd__o21ai_2 _3429_ (.A1(_2534_),
    .A2(_2533_),
    .B1(_2518_),
    .Y(_2589_));
 sky130_fd_sc_hd__nand3_1 _3430_ (.A(_2531_),
    .B(_2522_),
    .C(_2530_),
    .Y(_2590_));
 sky130_fd_sc_hd__a21o_1 _3431_ (.A1(_2531_),
    .A2(_2530_),
    .B1(_2522_),
    .X(_2591_));
 sky130_fd_sc_hd__xor2_1 _3432_ (.A(_2546_),
    .B(_2548_),
    .X(_2592_));
 sky130_fd_sc_hd__or3_1 _3433_ (.A(_2528_),
    .B(_2525_),
    .C(_2527_),
    .X(_2593_));
 sky130_fd_sc_hd__o21ai_1 _3434_ (.A1(_2528_),
    .A2(_2527_),
    .B1(_2525_),
    .Y(_2594_));
 sky130_fd_sc_hd__nand2_1 _3435_ (.A(_0960_),
    .B(_2438_),
    .Y(_2595_));
 sky130_fd_sc_hd__a22oi_2 _3436_ (.A1(_2496_),
    .A2(_0905_),
    .B1(_2238_),
    .B2(_2470_),
    .Y(_2596_));
 sky130_fd_sc_hd__and4_1 _3437_ (.A(\B[1][0] ),
    .B(\B[1][1] ),
    .C(\A[2][3] ),
    .D(\A[2][4] ),
    .X(_2597_));
 sky130_fd_sc_hd__o21bai_1 _3438_ (.A1(_2595_),
    .A2(_2596_),
    .B1_N(_2597_),
    .Y(_2598_));
 sky130_fd_sc_hd__a21o_1 _3439_ (.A1(_2593_),
    .A2(_2594_),
    .B1(_2598_),
    .X(_2599_));
 sky130_fd_sc_hd__nand3_1 _3440_ (.A(_2593_),
    .B(_2594_),
    .C(_2598_),
    .Y(_2600_));
 sky130_fd_sc_hd__a21bo_1 _3441_ (.A1(_2592_),
    .A2(_2599_),
    .B1_N(_2600_),
    .X(_2601_));
 sky130_fd_sc_hd__and3_1 _3442_ (.A(_2590_),
    .B(_2591_),
    .C(_2601_),
    .X(_2602_));
 sky130_fd_sc_hd__nand3_1 _3443_ (.A(_2590_),
    .B(_2591_),
    .C(_2601_),
    .Y(_2603_));
 sky130_fd_sc_hd__nor3_1 _3444_ (.A(_2545_),
    .B(_2549_),
    .C(_2553_),
    .Y(_2604_));
 sky130_fd_sc_hd__nor2_1 _3445_ (.A(_2554_),
    .B(_2604_),
    .Y(_2605_));
 sky130_fd_sc_hd__a21o_1 _3446_ (.A1(_2590_),
    .A2(_2591_),
    .B1(_2601_),
    .X(_2606_));
 sky130_fd_sc_hd__and3_1 _3447_ (.A(_2603_),
    .B(_2605_),
    .C(_2606_),
    .X(_2607_));
 sky130_fd_sc_hd__a211o_1 _3448_ (.A1(_2588_),
    .A2(_2589_),
    .B1(_2602_),
    .C1(_2607_),
    .X(_2608_));
 sky130_fd_sc_hd__o211ai_4 _3449_ (.A1(_2602_),
    .A2(_2607_),
    .B1(_2588_),
    .C1(_2589_),
    .Y(_2609_));
 sky130_fd_sc_hd__a21boi_1 _3450_ (.A1(_2587_),
    .A2(_2608_),
    .B1_N(_2609_),
    .Y(_2610_));
 sky130_fd_sc_hd__xnor2_1 _3451_ (.A(_2585_),
    .B(_2610_),
    .Y(_2611_));
 sky130_fd_sc_hd__nor2_1 _3452_ (.A(_2585_),
    .B(_2610_),
    .Y(_2612_));
 sky130_fd_sc_hd__o21ba_1 _3453_ (.A1(_2584_),
    .A2(_2611_),
    .B1_N(_2612_),
    .X(_2613_));
 sky130_fd_sc_hd__xnor2_1 _3454_ (.A(_2582_),
    .B(_2613_),
    .Y(_2614_));
 sky130_fd_sc_hd__and2b_1 _3455_ (.A_N(_2613_),
    .B(_2582_),
    .X(_2615_));
 sky130_fd_sc_hd__a21oi_1 _3456_ (.A1(_2581_),
    .A2(_2614_),
    .B1(_2615_),
    .Y(_2616_));
 sky130_fd_sc_hd__xor2_2 _3457_ (.A(_2543_),
    .B(_2616_),
    .X(_2617_));
 sky130_fd_sc_hd__and4_1 _3458_ (.A(_1312_),
    .B(_2568_),
    .C(_1598_),
    .D(_1334_),
    .X(_2618_));
 sky130_fd_sc_hd__and4_1 _3459_ (.A(\A[3][1] ),
    .B(_1136_),
    .C(_2559_),
    .D(_1103_),
    .X(_2619_));
 sky130_fd_sc_hd__a22oi_1 _3460_ (.A1(_1235_),
    .A2(_0707_),
    .B1(_1806_),
    .B2(_1598_),
    .Y(_2620_));
 sky130_fd_sc_hd__and4bb_1 _3461_ (.A_N(_2619_),
    .B_N(_2620_),
    .C(_2568_),
    .D(_2347_),
    .X(_2621_));
 sky130_fd_sc_hd__nor2_1 _3462_ (.A(_2619_),
    .B(_2621_),
    .Y(_2622_));
 sky130_fd_sc_hd__nand2_1 _3463_ (.A(_1609_),
    .B(_2347_),
    .Y(_2623_));
 sky130_fd_sc_hd__and4_1 _3464_ (.A(_1092_),
    .B(_2559_),
    .C(_1257_),
    .D(\A[3][3] ),
    .X(_2624_));
 sky130_fd_sc_hd__a22o_1 _3465_ (.A1(_2559_),
    .A2(_1257_),
    .B1(_1323_),
    .B2(_1136_),
    .X(_2625_));
 sky130_fd_sc_hd__and2b_1 _3466_ (.A_N(_2624_),
    .B(_2625_),
    .X(_2626_));
 sky130_fd_sc_hd__xnor2_1 _3467_ (.A(_2623_),
    .B(_2626_),
    .Y(_2627_));
 sky130_fd_sc_hd__and2b_1 _3468_ (.A_N(_2622_),
    .B(_2627_),
    .X(_2628_));
 sky130_fd_sc_hd__buf_2 _3469_ (.A(_2568_),
    .X(_2629_));
 sky130_fd_sc_hd__buf_4 _3470_ (.A(_1543_),
    .X(_2630_));
 sky130_fd_sc_hd__xnor2_1 _3471_ (.A(_2627_),
    .B(_2622_),
    .Y(_2631_));
 sky130_fd_sc_hd__and3_1 _3472_ (.A(_2629_),
    .B(_2630_),
    .C(_2631_),
    .X(_2632_));
 sky130_fd_sc_hd__a22oi_1 _3473_ (.A1(_1521_),
    .A2(_2568_),
    .B1(_1609_),
    .B2(_1543_),
    .Y(_2633_));
 sky130_fd_sc_hd__or2_1 _3474_ (.A(_2618_),
    .B(_2633_),
    .X(_2634_));
 sky130_fd_sc_hd__or3_1 _3475_ (.A(_2562_),
    .B(_2560_),
    .C(_2561_),
    .X(_2635_));
 sky130_fd_sc_hd__o21ai_1 _3476_ (.A1(_2562_),
    .A2(_2561_),
    .B1(_2560_),
    .Y(_2636_));
 sky130_fd_sc_hd__a31o_1 _3477_ (.A1(_1598_),
    .A2(_1202_),
    .A3(_2625_),
    .B1(_2624_),
    .X(_2637_));
 sky130_fd_sc_hd__and3_1 _3478_ (.A(_2635_),
    .B(_2636_),
    .C(_2637_),
    .X(_2638_));
 sky130_fd_sc_hd__a21oi_1 _3479_ (.A1(_2635_),
    .A2(_2636_),
    .B1(_2637_),
    .Y(_2639_));
 sky130_fd_sc_hd__nor2_1 _3480_ (.A(_2638_),
    .B(_2639_),
    .Y(_2640_));
 sky130_fd_sc_hd__xnor2_1 _3481_ (.A(_2634_),
    .B(_2640_),
    .Y(_2641_));
 sky130_fd_sc_hd__o21a_1 _3482_ (.A1(_2628_),
    .A2(_2632_),
    .B1(_2641_),
    .X(_2642_));
 sky130_fd_sc_hd__and2_1 _3483_ (.A(_2618_),
    .B(_2642_),
    .X(_2643_));
 sky130_fd_sc_hd__or3_1 _3484_ (.A(_2597_),
    .B(_2595_),
    .C(_2596_),
    .X(_2644_));
 sky130_fd_sc_hd__o21ai_1 _3485_ (.A1(_2597_),
    .A2(_2596_),
    .B1(_2595_),
    .Y(_2645_));
 sky130_fd_sc_hd__nand2_1 _3486_ (.A(_0817_),
    .B(_2438_),
    .Y(_2646_));
 sky130_fd_sc_hd__a22oi_2 _3487_ (.A1(_2496_),
    .A2(_0960_),
    .B1(_1004_),
    .B2(_2470_),
    .Y(_2647_));
 sky130_fd_sc_hd__and4_1 _3488_ (.A(\B[1][0] ),
    .B(\B[1][1] ),
    .C(_0960_),
    .D(_0905_),
    .X(_2648_));
 sky130_fd_sc_hd__o21bai_1 _3489_ (.A1(_2646_),
    .A2(_2647_),
    .B1_N(_2648_),
    .Y(_2649_));
 sky130_fd_sc_hd__nand3_1 _3490_ (.A(_2644_),
    .B(_2645_),
    .C(_2649_),
    .Y(_2650_));
 sky130_fd_sc_hd__and4_1 _3491_ (.A(_0762_),
    .B(_0817_),
    .C(_0927_),
    .D(_0949_),
    .X(_2651_));
 sky130_fd_sc_hd__a22oi_1 _3492_ (.A1(_0883_),
    .A2(_2440_),
    .B1(_0949_),
    .B2(_0773_),
    .Y(_2652_));
 sky130_fd_sc_hd__nor2_1 _3493_ (.A(_2651_),
    .B(_2652_),
    .Y(_2653_));
 sky130_fd_sc_hd__a21o_1 _3494_ (.A1(_2644_),
    .A2(_2645_),
    .B1(_2649_),
    .X(_2654_));
 sky130_fd_sc_hd__nand3_1 _3495_ (.A(_2650_),
    .B(_2653_),
    .C(_2654_),
    .Y(_2655_));
 sky130_fd_sc_hd__a21o_1 _3496_ (.A1(_2650_),
    .A2(_2654_),
    .B1(_2653_),
    .X(_2656_));
 sky130_fd_sc_hd__nand2_1 _3497_ (.A(_2550_),
    .B(_2440_),
    .Y(_2657_));
 sky130_fd_sc_hd__or3_1 _3498_ (.A(_2648_),
    .B(_2646_),
    .C(_2647_),
    .X(_2658_));
 sky130_fd_sc_hd__o21ai_1 _3499_ (.A1(_2648_),
    .A2(_2647_),
    .B1(_2646_),
    .Y(_2659_));
 sky130_fd_sc_hd__a22o_1 _3500_ (.A1(_0872_),
    .A2(_2437_),
    .B1(_0960_),
    .B2(_2468_),
    .X(_2660_));
 sky130_fd_sc_hd__and4_1 _3501_ (.A(_2468_),
    .B(_0872_),
    .C(_2496_),
    .D(_0960_),
    .X(_2661_));
 sky130_fd_sc_hd__a31o_1 _3502_ (.A1(_0762_),
    .A2(_2432_),
    .A3(_2660_),
    .B1(_2661_),
    .X(_2662_));
 sky130_fd_sc_hd__a21oi_2 _3503_ (.A1(_2658_),
    .A2(_2659_),
    .B1(_2662_),
    .Y(_2663_));
 sky130_fd_sc_hd__and3_1 _3504_ (.A(_2658_),
    .B(_2659_),
    .C(_2662_),
    .X(_2664_));
 sky130_fd_sc_hd__o21bai_2 _3505_ (.A1(_2657_),
    .A2(_2663_),
    .B1_N(_2664_),
    .Y(_2665_));
 sky130_fd_sc_hd__nand3_4 _3506_ (.A(_2655_),
    .B(_2656_),
    .C(_2665_),
    .Y(_2666_));
 sky130_fd_sc_hd__buf_4 _3507_ (.A(_0784_),
    .X(_2667_));
 sky130_fd_sc_hd__buf_4 _3508_ (.A(_1213_),
    .X(_2668_));
 sky130_fd_sc_hd__a21o_1 _3509_ (.A1(_2655_),
    .A2(_2656_),
    .B1(_2665_),
    .X(_2669_));
 sky130_fd_sc_hd__nand4_4 _3510_ (.A(_2667_),
    .B(_2668_),
    .C(_2666_),
    .D(_2669_),
    .Y(_2670_));
 sky130_fd_sc_hd__nand3_1 _3511_ (.A(_2600_),
    .B(_2592_),
    .C(_2599_),
    .Y(_2671_));
 sky130_fd_sc_hd__a21o_1 _3512_ (.A1(_2600_),
    .A2(_2599_),
    .B1(_2592_),
    .X(_2672_));
 sky130_fd_sc_hd__a21bo_1 _3513_ (.A1(_2653_),
    .A2(_2654_),
    .B1_N(_2650_),
    .X(_2673_));
 sky130_fd_sc_hd__and3_2 _3514_ (.A(_2671_),
    .B(_2672_),
    .C(_2673_),
    .X(_2674_));
 sky130_fd_sc_hd__and3_1 _3515_ (.A(_1740_),
    .B(_0784_),
    .C(_2651_),
    .X(_2675_));
 sky130_fd_sc_hd__clkbuf_4 _3516_ (.A(_1740_),
    .X(_2676_));
 sky130_fd_sc_hd__a21oi_1 _3517_ (.A1(_2676_),
    .A2(_0784_),
    .B1(_2651_),
    .Y(_2677_));
 sky130_fd_sc_hd__or2_1 _3518_ (.A(_2675_),
    .B(_2677_),
    .X(_2678_));
 sky130_fd_sc_hd__a21oi_2 _3519_ (.A1(_2671_),
    .A2(_2672_),
    .B1(_2673_),
    .Y(_2679_));
 sky130_fd_sc_hd__nor3_4 _3520_ (.A(_2674_),
    .B(_2678_),
    .C(_2679_),
    .Y(_2680_));
 sky130_fd_sc_hd__o21a_1 _3521_ (.A1(_2674_),
    .A2(_2679_),
    .B1(_2678_),
    .X(_2681_));
 sky130_fd_sc_hd__a211oi_4 _3522_ (.A1(_2666_),
    .A2(_2670_),
    .B1(_2680_),
    .C1(_2681_),
    .Y(_2682_));
 sky130_fd_sc_hd__inv_2 _3523_ (.A(_2682_),
    .Y(_2683_));
 sky130_fd_sc_hd__o211a_1 _3524_ (.A1(_2680_),
    .A2(_2681_),
    .B1(_2666_),
    .C1(_2670_),
    .X(_2684_));
 sky130_fd_sc_hd__nor3_1 _3525_ (.A(_2628_),
    .B(_2632_),
    .C(_2641_),
    .Y(_2685_));
 sky130_fd_sc_hd__nor2_1 _3526_ (.A(_2642_),
    .B(_2685_),
    .Y(_2686_));
 sky130_fd_sc_hd__or3b_4 _3527_ (.A(_2682_),
    .B(_2684_),
    .C_N(_2686_),
    .X(_2687_));
 sky130_fd_sc_hd__nand3_1 _3528_ (.A(_2603_),
    .B(_2605_),
    .C(_2606_),
    .Y(_2688_));
 sky130_fd_sc_hd__a21o_1 _3529_ (.A1(_2603_),
    .A2(_2606_),
    .B1(_2605_),
    .X(_2689_));
 sky130_fd_sc_hd__o211a_2 _3530_ (.A1(_2674_),
    .A2(_2680_),
    .B1(_2688_),
    .C1(_2689_),
    .X(_2690_));
 sky130_fd_sc_hd__o21ba_1 _3531_ (.A1(_2634_),
    .A2(_2639_),
    .B1_N(_2638_),
    .X(_2691_));
 sky130_fd_sc_hd__inv_2 _3532_ (.A(_2691_),
    .Y(_2692_));
 sky130_fd_sc_hd__a21o_1 _3533_ (.A1(_2564_),
    .A2(_2571_),
    .B1(_2570_),
    .X(_2693_));
 sky130_fd_sc_hd__nand3_1 _3534_ (.A(_2572_),
    .B(_2675_),
    .C(_2693_),
    .Y(_2694_));
 sky130_fd_sc_hd__a21o_1 _3535_ (.A1(_2572_),
    .A2(_2693_),
    .B1(_2675_),
    .X(_2695_));
 sky130_fd_sc_hd__and3_1 _3536_ (.A(_2692_),
    .B(_2694_),
    .C(_2695_),
    .X(_2696_));
 sky130_fd_sc_hd__a21oi_1 _3537_ (.A1(_2694_),
    .A2(_2695_),
    .B1(_2692_),
    .Y(_2697_));
 sky130_fd_sc_hd__or2_1 _3538_ (.A(_2696_),
    .B(_2697_),
    .X(_2698_));
 sky130_fd_sc_hd__a211oi_4 _3539_ (.A1(_2688_),
    .A2(_2689_),
    .B1(_2674_),
    .C1(_2680_),
    .Y(_2699_));
 sky130_fd_sc_hd__nor3_2 _3540_ (.A(_2690_),
    .B(_2698_),
    .C(_2699_),
    .Y(_2700_));
 sky130_fd_sc_hd__o21a_1 _3541_ (.A1(_2690_),
    .A2(_2699_),
    .B1(_2698_),
    .X(_2701_));
 sky130_fd_sc_hd__a211oi_4 _3542_ (.A1(_2683_),
    .A2(_2687_),
    .B1(_2700_),
    .C1(_2701_),
    .Y(_2702_));
 sky130_fd_sc_hd__nor2_1 _3543_ (.A(_2618_),
    .B(_2642_),
    .Y(_2703_));
 sky130_fd_sc_hd__or2_1 _3544_ (.A(_2643_),
    .B(_2703_),
    .X(_2704_));
 sky130_fd_sc_hd__o211a_1 _3545_ (.A1(_2700_),
    .A2(_2701_),
    .B1(_2683_),
    .C1(_2687_),
    .X(_2705_));
 sky130_fd_sc_hd__nor3_2 _3546_ (.A(_2702_),
    .B(_2704_),
    .C(_2705_),
    .Y(_2706_));
 sky130_fd_sc_hd__inv_2 _3547_ (.A(_2690_),
    .Y(_2707_));
 sky130_fd_sc_hd__or3_1 _3548_ (.A(_2690_),
    .B(_2698_),
    .C(_2699_),
    .X(_2708_));
 sky130_fd_sc_hd__and3_1 _3549_ (.A(_2609_),
    .B(_2587_),
    .C(_2608_),
    .X(_2709_));
 sky130_fd_sc_hd__a21oi_1 _3550_ (.A1(_2609_),
    .A2(_2608_),
    .B1(_2587_),
    .Y(_2710_));
 sky130_fd_sc_hd__a211o_1 _3551_ (.A1(_2707_),
    .A2(_2708_),
    .B1(_2709_),
    .C1(_2710_),
    .X(_2711_));
 sky130_fd_sc_hd__and3_1 _3552_ (.A(_2572_),
    .B(_2675_),
    .C(_2693_),
    .X(_2712_));
 sky130_fd_sc_hd__o21ba_1 _3553_ (.A1(_2565_),
    .A2(_2569_),
    .B1_N(_2566_),
    .X(_2713_));
 sky130_fd_sc_hd__o21ba_1 _3554_ (.A1(_2712_),
    .A2(_2696_),
    .B1_N(_2713_),
    .X(_2714_));
 sky130_fd_sc_hd__or3b_1 _3555_ (.A(_2712_),
    .B(_2696_),
    .C_N(_2713_),
    .X(_2715_));
 sky130_fd_sc_hd__and2b_1 _3556_ (.A_N(_2714_),
    .B(_2715_),
    .X(_2716_));
 sky130_fd_sc_hd__clkbuf_4 _3557_ (.A(_2629_),
    .X(_2717_));
 sky130_fd_sc_hd__nand2_1 _3558_ (.A(_0674_),
    .B(_2717_),
    .Y(_2718_));
 sky130_fd_sc_hd__xnor2_1 _3559_ (.A(_2716_),
    .B(_2718_),
    .Y(_2719_));
 sky130_fd_sc_hd__o211ai_2 _3560_ (.A1(_2709_),
    .A2(_2710_),
    .B1(_2707_),
    .C1(_2708_),
    .Y(_2720_));
 sky130_fd_sc_hd__nand3_1 _3561_ (.A(_2711_),
    .B(_2719_),
    .C(_2720_),
    .Y(_2721_));
 sky130_fd_sc_hd__a21o_1 _3562_ (.A1(_2711_),
    .A2(_2720_),
    .B1(_2719_),
    .X(_2722_));
 sky130_fd_sc_hd__o211ai_2 _3563_ (.A1(_2702_),
    .A2(_2706_),
    .B1(_2721_),
    .C1(_2722_),
    .Y(_2723_));
 sky130_fd_sc_hd__a211o_1 _3564_ (.A1(_2721_),
    .A2(_2722_),
    .B1(_2702_),
    .C1(_2706_),
    .X(_2724_));
 sky130_fd_sc_hd__and3_1 _3565_ (.A(_2643_),
    .B(_2723_),
    .C(_2724_),
    .X(_2725_));
 sky130_fd_sc_hd__a21oi_1 _3566_ (.A1(_2723_),
    .A2(_2724_),
    .B1(_2643_),
    .Y(_2726_));
 sky130_fd_sc_hd__a22o_1 _3567_ (.A1(_2667_),
    .A2(_2668_),
    .B1(_2666_),
    .B2(_2669_),
    .X(_2727_));
 sky130_fd_sc_hd__and2_1 _3568_ (.A(_2667_),
    .B(_1532_),
    .X(_2728_));
 sky130_fd_sc_hd__or3_1 _3569_ (.A(_2657_),
    .B(_2664_),
    .C(_2663_),
    .X(_2729_));
 sky130_fd_sc_hd__o21ai_2 _3570_ (.A1(_2664_),
    .A2(_2663_),
    .B1(_2657_),
    .Y(_2730_));
 sky130_fd_sc_hd__nand2_1 _3571_ (.A(_0773_),
    .B(_2432_),
    .Y(_2731_));
 sky130_fd_sc_hd__and2b_1 _3572_ (.A_N(_2661_),
    .B(_2660_),
    .X(_2732_));
 sky130_fd_sc_hd__xnor2_2 _3573_ (.A(_2731_),
    .B(_2732_),
    .Y(_2733_));
 sky130_fd_sc_hd__and4_1 _3574_ (.A(_2471_),
    .B(_0773_),
    .C(_0883_),
    .D(_2433_),
    .X(_2734_));
 sky130_fd_sc_hd__and2_1 _3575_ (.A(_2733_),
    .B(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__a21o_1 _3576_ (.A1(_2729_),
    .A2(_2730_),
    .B1(_2735_),
    .X(_2736_));
 sky130_fd_sc_hd__nand3_1 _3577_ (.A(_2729_),
    .B(_2730_),
    .C(_2735_),
    .Y(_2737_));
 sky130_fd_sc_hd__a21bo_1 _3578_ (.A1(_2728_),
    .A2(_2736_),
    .B1_N(_2737_),
    .X(_2738_));
 sky130_fd_sc_hd__and3_2 _3579_ (.A(_2670_),
    .B(_2727_),
    .C(_2738_),
    .X(_2739_));
 sky130_fd_sc_hd__nand2_1 _3580_ (.A(_2629_),
    .B(_2630_),
    .Y(_2740_));
 sky130_fd_sc_hd__xnor2_1 _3581_ (.A(_2740_),
    .B(_2631_),
    .Y(_2741_));
 sky130_fd_sc_hd__o2bb2a_1 _3582_ (.A1_N(_2568_),
    .A2_N(_2347_),
    .B1(_2619_),
    .B2(_2620_),
    .X(_2742_));
 sky130_fd_sc_hd__nor2_1 _3583_ (.A(_2621_),
    .B(_2742_),
    .Y(_2743_));
 sky130_fd_sc_hd__and4_1 _3584_ (.A(_2629_),
    .B(_1609_),
    .C(_1235_),
    .D(_1806_),
    .X(_2744_));
 sky130_fd_sc_hd__and2_1 _3585_ (.A(_2743_),
    .B(_2744_),
    .X(_2745_));
 sky130_fd_sc_hd__and2_1 _3586_ (.A(_2741_),
    .B(_2745_),
    .X(_2746_));
 sky130_fd_sc_hd__nor2_1 _3587_ (.A(_2741_),
    .B(_2745_),
    .Y(_2747_));
 sky130_fd_sc_hd__or2_1 _3588_ (.A(_2746_),
    .B(_2747_),
    .X(_2748_));
 sky130_fd_sc_hd__a21oi_1 _3589_ (.A1(_2670_),
    .A2(_2727_),
    .B1(_2738_),
    .Y(_2749_));
 sky130_fd_sc_hd__nor3_1 _3590_ (.A(_2739_),
    .B(_2748_),
    .C(_2749_),
    .Y(_2750_));
 sky130_fd_sc_hd__o21bai_2 _3591_ (.A1(_2682_),
    .A2(_2684_),
    .B1_N(_2686_),
    .Y(_2751_));
 sky130_fd_sc_hd__o211ai_4 _3592_ (.A1(_2739_),
    .A2(_2750_),
    .B1(_2687_),
    .C1(_2751_),
    .Y(_2752_));
 sky130_fd_sc_hd__a211o_1 _3593_ (.A1(_2687_),
    .A2(_2751_),
    .B1(_2739_),
    .C1(_2750_),
    .X(_2753_));
 sky130_fd_sc_hd__nand3_2 _3594_ (.A(_2746_),
    .B(_2752_),
    .C(_2753_),
    .Y(_2754_));
 sky130_fd_sc_hd__o21a_1 _3595_ (.A1(_2702_),
    .A2(_2705_),
    .B1(_2704_),
    .X(_2755_));
 sky130_fd_sc_hd__a211oi_2 _3596_ (.A1(_2752_),
    .A2(_2754_),
    .B1(_2755_),
    .C1(_2706_),
    .Y(_2756_));
 sky130_fd_sc_hd__o211a_1 _3597_ (.A1(_2706_),
    .A2(_2755_),
    .B1(_2754_),
    .C1(_2752_),
    .X(_2757_));
 sky130_fd_sc_hd__a21o_1 _3598_ (.A1(_2752_),
    .A2(_2753_),
    .B1(_2746_),
    .X(_2758_));
 sky130_fd_sc_hd__and2_1 _3599_ (.A(_2754_),
    .B(_2758_),
    .X(_2759_));
 sky130_fd_sc_hd__or3_1 _3600_ (.A(_2739_),
    .B(_2748_),
    .C(_2749_),
    .X(_2760_));
 sky130_fd_sc_hd__o21ai_1 _3601_ (.A1(_2739_),
    .A2(_2749_),
    .B1(_2748_),
    .Y(_2761_));
 sky130_fd_sc_hd__nand3_1 _3602_ (.A(_2737_),
    .B(_2728_),
    .C(_2736_),
    .Y(_2762_));
 sky130_fd_sc_hd__a21o_1 _3603_ (.A1(_2737_),
    .A2(_2736_),
    .B1(_2728_),
    .X(_2763_));
 sky130_fd_sc_hd__inv_2 _3604_ (.A(_2734_),
    .Y(_2764_));
 sky130_fd_sc_hd__xnor2_1 _3605_ (.A(_2733_),
    .B(_2764_),
    .Y(_2765_));
 sky130_fd_sc_hd__and3_1 _3606_ (.A(_2667_),
    .B(_0718_),
    .C(_2765_),
    .X(_2766_));
 sky130_fd_sc_hd__a21o_1 _3607_ (.A1(_2762_),
    .A2(_2763_),
    .B1(_2766_),
    .X(_2767_));
 sky130_fd_sc_hd__nor2_1 _3608_ (.A(_2743_),
    .B(_2744_),
    .Y(_2768_));
 sky130_fd_sc_hd__nor2_1 _3609_ (.A(_2745_),
    .B(_2768_),
    .Y(_2769_));
 sky130_fd_sc_hd__nand3_1 _3610_ (.A(_2762_),
    .B(_2763_),
    .C(_2766_),
    .Y(_2770_));
 sky130_fd_sc_hd__a21bo_1 _3611_ (.A1(_2767_),
    .A2(_2769_),
    .B1_N(_2770_),
    .X(_2771_));
 sky130_fd_sc_hd__and3_1 _3612_ (.A(_2760_),
    .B(_2761_),
    .C(_2771_),
    .X(_2772_));
 sky130_fd_sc_hd__or4bb_2 _3613_ (.A(_2756_),
    .B(_2757_),
    .C_N(_2759_),
    .D_N(_2772_),
    .X(_2773_));
 sky130_fd_sc_hd__and2b_1 _3614_ (.A_N(_2756_),
    .B(_2773_),
    .X(_2774_));
 sky130_fd_sc_hd__a21o_1 _3615_ (.A1(_2760_),
    .A2(_2761_),
    .B1(_2771_),
    .X(_2775_));
 sky130_fd_sc_hd__nand2_1 _3616_ (.A(_2770_),
    .B(_2767_),
    .Y(_2776_));
 sky130_fd_sc_hd__xnor2_1 _3617_ (.A(_2776_),
    .B(_2769_),
    .Y(_2777_));
 sky130_fd_sc_hd__clkbuf_4 _3618_ (.A(_2667_),
    .X(_2778_));
 sky130_fd_sc_hd__a21oi_1 _3619_ (.A1(_2778_),
    .A2(_0718_),
    .B1(_2765_),
    .Y(_2779_));
 sky130_fd_sc_hd__nor2_1 _3620_ (.A(_2766_),
    .B(_2779_),
    .Y(_2780_));
 sky130_fd_sc_hd__a22o_1 _3621_ (.A1(_2471_),
    .A2(_0883_),
    .B1(_2433_),
    .B2(_2550_),
    .X(_2781_));
 sky130_fd_sc_hd__and4_1 _3622_ (.A(_2778_),
    .B(_2544_),
    .C(_2764_),
    .D(_2781_),
    .X(_2782_));
 sky130_fd_sc_hd__xnor2_1 _3623_ (.A(_2780_),
    .B(_2782_),
    .Y(_2783_));
 sky130_fd_sc_hd__a22oi_1 _3624_ (.A1(_2544_),
    .A2(_1235_),
    .B1(_1806_),
    .B2(_2629_),
    .Y(_2784_));
 sky130_fd_sc_hd__or2_1 _3625_ (.A(_2744_),
    .B(_2784_),
    .X(_2785_));
 sky130_fd_sc_hd__nor2_1 _3626_ (.A(_2783_),
    .B(_2785_),
    .Y(_2786_));
 sky130_fd_sc_hd__a21o_1 _3627_ (.A1(_2780_),
    .A2(_2782_),
    .B1(_2786_),
    .X(_2787_));
 sky130_fd_sc_hd__and4b_1 _3628_ (.A_N(_2772_),
    .B(_2775_),
    .C(_2777_),
    .D(_2787_),
    .X(_2788_));
 sky130_fd_sc_hd__and3_1 _3629_ (.A(_2754_),
    .B(_2788_),
    .C(_2758_),
    .X(_2789_));
 sky130_fd_sc_hd__and2b_1 _3630_ (.A_N(_2772_),
    .B(_2775_),
    .X(_2790_));
 sky130_fd_sc_hd__xor2_1 _3631_ (.A(_2777_),
    .B(_2787_),
    .X(_2791_));
 sky130_fd_sc_hd__and2_1 _3632_ (.A(_2783_),
    .B(_2785_),
    .X(_2792_));
 sky130_fd_sc_hd__nor2_1 _3633_ (.A(_2786_),
    .B(_2792_),
    .Y(_2793_));
 sky130_fd_sc_hd__a22oi_1 _3634_ (.A1(_2778_),
    .A2(_2544_),
    .B1(_2764_),
    .B2(_2781_),
    .Y(_2794_));
 sky130_fd_sc_hd__nor2_1 _3635_ (.A(_2782_),
    .B(_2794_),
    .Y(_2795_));
 sky130_fd_sc_hd__and4_1 _3636_ (.A(_2471_),
    .B(_2550_),
    .C(_2629_),
    .D(_2778_),
    .X(_2796_));
 sky130_fd_sc_hd__nand2_1 _3637_ (.A(_2717_),
    .B(_1235_),
    .Y(_2797_));
 sky130_fd_sc_hd__xnor2_1 _3638_ (.A(_2795_),
    .B(_2796_),
    .Y(_2798_));
 sky130_fd_sc_hd__nor2_1 _3639_ (.A(_2797_),
    .B(_2798_),
    .Y(_2799_));
 sky130_fd_sc_hd__a21o_1 _3640_ (.A1(_2795_),
    .A2(_2796_),
    .B1(_2799_),
    .X(_2800_));
 sky130_fd_sc_hd__and2_1 _3641_ (.A(_2793_),
    .B(_2800_),
    .X(_2801_));
 sky130_fd_sc_hd__and3_1 _3642_ (.A(_2790_),
    .B(_2791_),
    .C(_2801_),
    .X(_2802_));
 sky130_fd_sc_hd__a211o_1 _3643_ (.A1(_2754_),
    .A2(_2758_),
    .B1(_2788_),
    .C1(_2772_),
    .X(_2803_));
 sky130_fd_sc_hd__o211ai_1 _3644_ (.A1(_2772_),
    .A2(_2788_),
    .B1(_2758_),
    .C1(_2754_),
    .Y(_2804_));
 sky130_fd_sc_hd__and3_1 _3645_ (.A(_2802_),
    .B(_2803_),
    .C(_2804_),
    .X(_2805_));
 sky130_fd_sc_hd__a2bb2o_1 _3646_ (.A1_N(_2756_),
    .A2_N(_2757_),
    .B1(_2759_),
    .B2(_2772_),
    .X(_2806_));
 sky130_fd_sc_hd__o211ai_4 _3647_ (.A1(_2789_),
    .A2(_2805_),
    .B1(_2773_),
    .C1(_2806_),
    .Y(_2807_));
 sky130_fd_sc_hd__nand3_1 _3648_ (.A(_2643_),
    .B(_2723_),
    .C(_2724_),
    .Y(_2808_));
 sky130_fd_sc_hd__a21o_1 _3649_ (.A1(_2723_),
    .A2(_2724_),
    .B1(_2643_),
    .X(_2809_));
 sky130_fd_sc_hd__a21oi_2 _3650_ (.A1(_2808_),
    .A2(_2809_),
    .B1(_2756_),
    .Y(_2810_));
 sky130_fd_sc_hd__o32ai_4 _3651_ (.A1(_2725_),
    .A2(_2726_),
    .A3(_2774_),
    .B1(_2807_),
    .B2(_2810_),
    .Y(_2811_));
 sky130_fd_sc_hd__a31o_1 _3652_ (.A1(_0685_),
    .A2(_2717_),
    .A3(_2716_),
    .B1(_2714_),
    .X(_2812_));
 sky130_fd_sc_hd__xnor2_2 _3653_ (.A(_2584_),
    .B(_2611_),
    .Y(_2813_));
 sky130_fd_sc_hd__a21bo_1 _3654_ (.A1(_2719_),
    .A2(_2720_),
    .B1_N(_2711_),
    .X(_2814_));
 sky130_fd_sc_hd__xnor2_2 _3655_ (.A(_2813_),
    .B(_2814_),
    .Y(_2815_));
 sky130_fd_sc_hd__xor2_2 _3656_ (.A(_2812_),
    .B(_2815_),
    .X(_2816_));
 sky130_fd_sc_hd__a21bo_1 _3657_ (.A1(_2643_),
    .A2(_2724_),
    .B1_N(_2723_),
    .X(_2817_));
 sky130_fd_sc_hd__xor2_1 _3658_ (.A(_2816_),
    .B(_2817_),
    .X(_2818_));
 sky130_fd_sc_hd__xnor2_2 _3659_ (.A(_2581_),
    .B(_2614_),
    .Y(_2819_));
 sky130_fd_sc_hd__or2b_1 _3660_ (.A(_2813_),
    .B_N(_2814_),
    .X(_2820_));
 sky130_fd_sc_hd__a21boi_2 _3661_ (.A1(_2812_),
    .A2(_2815_),
    .B1_N(_2820_),
    .Y(_2821_));
 sky130_fd_sc_hd__xor2_2 _3662_ (.A(_2819_),
    .B(_2821_),
    .X(_2822_));
 sky130_fd_sc_hd__a2bb2o_1 _3663_ (.A1_N(_2819_),
    .A2_N(_2821_),
    .B1(_2816_),
    .B2(_2817_),
    .X(_2823_));
 sky130_fd_sc_hd__a21boi_1 _3664_ (.A1(_2819_),
    .A2(_2821_),
    .B1_N(_2823_),
    .Y(_2824_));
 sky130_fd_sc_hd__a31o_1 _3665_ (.A1(_2811_),
    .A2(_2818_),
    .A3(_2822_),
    .B1(_2824_),
    .X(_2825_));
 sky130_fd_sc_hd__or2_1 _3666_ (.A(_2543_),
    .B(_2616_),
    .X(_2826_));
 sky130_fd_sc_hd__a21bo_1 _3667_ (.A1(_2617_),
    .A2(_2825_),
    .B1_N(_2826_),
    .X(_2827_));
 sky130_fd_sc_hd__nor2_1 _3668_ (.A(_2509_),
    .B(_2541_),
    .Y(_2828_));
 sky130_fd_sc_hd__a21oi_2 _3669_ (.A1(_1729_),
    .A2(_2542_),
    .B1(_2828_),
    .Y(_2829_));
 sky130_fd_sc_hd__a31o_1 _3670_ (.A1(_0696_),
    .A2(_1532_),
    .A3(_2112_),
    .B1(_2090_),
    .X(_2830_));
 sky130_fd_sc_hd__nor2_1 _3671_ (.A(_2483_),
    .B(_2507_),
    .Y(_2831_));
 sky130_fd_sc_hd__a21o_1 _3672_ (.A1(_2133_),
    .A2(_2508_),
    .B1(_2831_),
    .X(_2832_));
 sky130_fd_sc_hd__clkbuf_4 _3673_ (.A(_1587_),
    .X(_2833_));
 sky130_fd_sc_hd__a32o_1 _3674_ (.A1(_2833_),
    .A2(_2668_),
    .A3(_2310_),
    .B1(_2300_),
    .B2(_2630_),
    .X(_2834_));
 sky130_fd_sc_hd__a21o_1 _3675_ (.A1(_2177_),
    .A2(_2373_),
    .B1(_2367_),
    .X(_2835_));
 sky130_fd_sc_hd__xor2_1 _3676_ (.A(_2834_),
    .B(_2835_),
    .X(_2836_));
 sky130_fd_sc_hd__and3_1 _3677_ (.A(\B[3][7] ),
    .B(_2668_),
    .C(_2836_),
    .X(_2837_));
 sky130_fd_sc_hd__a21oi_1 _3678_ (.A1(_0674_),
    .A2(_2668_),
    .B1(_2836_),
    .Y(_2838_));
 sky130_fd_sc_hd__nor2_1 _3679_ (.A(_2837_),
    .B(_2838_),
    .Y(_2839_));
 sky130_fd_sc_hd__and2_1 _3680_ (.A(_2460_),
    .B(_2481_),
    .X(_2840_));
 sky130_fd_sc_hd__a21oi_2 _3681_ (.A1(_2385_),
    .A2(_2482_),
    .B1(_2840_),
    .Y(_2841_));
 sky130_fd_sc_hd__a21oi_2 _3682_ (.A1(_2340_),
    .A2(_2354_),
    .B1(_2155_),
    .Y(_2842_));
 sky130_fd_sc_hd__and2b_1 _3683_ (.A_N(_2455_),
    .B(_2451_),
    .X(_2843_));
 sky130_fd_sc_hd__nand2_1 _3684_ (.A(_1587_),
    .B(_2676_),
    .Y(_2844_));
 sky130_fd_sc_hd__buf_2 _3685_ (.A(_0806_),
    .X(_2845_));
 sky130_fd_sc_hd__and2_1 _3686_ (.A(_1521_),
    .B(_0751_),
    .X(_2846_));
 sky130_fd_sc_hd__a21oi_1 _3687_ (.A1(_2845_),
    .A2(_2630_),
    .B1(_2846_),
    .Y(_2847_));
 sky130_fd_sc_hd__and3_1 _3688_ (.A(_0806_),
    .B(_2630_),
    .C(_2846_),
    .X(_2848_));
 sky130_fd_sc_hd__nor2_1 _3689_ (.A(_2847_),
    .B(_2848_),
    .Y(_2849_));
 sky130_fd_sc_hd__xnor2_1 _3690_ (.A(_2844_),
    .B(_2849_),
    .Y(_2850_));
 sky130_fd_sc_hd__o21a_1 _3691_ (.A1(_2843_),
    .A2(_2458_),
    .B1(_2850_),
    .X(_2851_));
 sky130_fd_sc_hd__nor3_1 _3692_ (.A(_2843_),
    .B(_2458_),
    .C(_2850_),
    .Y(_2852_));
 sky130_fd_sc_hd__nor2_1 _3693_ (.A(_2851_),
    .B(_2852_),
    .Y(_2853_));
 sky130_fd_sc_hd__xnor2_2 _3694_ (.A(_2842_),
    .B(_2853_),
    .Y(_2854_));
 sky130_fd_sc_hd__a21oi_2 _3695_ (.A1(_2449_),
    .A2(_2459_),
    .B1(_2448_),
    .Y(_2855_));
 sky130_fd_sc_hd__clkbuf_4 _3696_ (.A(_1904_),
    .X(_2856_));
 sky130_fd_sc_hd__nand2_2 _3697_ (.A(_2431_),
    .B(_2856_),
    .Y(_2857_));
 sky130_fd_sc_hd__buf_2 _3698_ (.A(_2405_),
    .X(_2858_));
 sky130_fd_sc_hd__clkbuf_4 _3699_ (.A(_2431_),
    .X(_2859_));
 sky130_fd_sc_hd__a22o_1 _3700_ (.A1(_2856_),
    .A2(_2858_),
    .B1(_0949_),
    .B2(_2859_),
    .X(_2860_));
 sky130_fd_sc_hd__o21ai_2 _3701_ (.A1(_2442_),
    .A2(_2857_),
    .B1(_2860_),
    .Y(_2861_));
 sky130_fd_sc_hd__clkbuf_4 _3702_ (.A(_1959_),
    .X(_2862_));
 sky130_fd_sc_hd__a22o_1 _3703_ (.A1(_0740_),
    .A2(_2445_),
    .B1(_2862_),
    .B2(_1915_),
    .X(_2863_));
 sky130_fd_sc_hd__nand2_1 _3704_ (.A(_2445_),
    .B(_1959_),
    .Y(_2864_));
 sky130_fd_sc_hd__or2_1 _3705_ (.A(_2453_),
    .B(_2864_),
    .X(_2865_));
 sky130_fd_sc_hd__nand2_1 _3706_ (.A(_2863_),
    .B(_2865_),
    .Y(_2866_));
 sky130_fd_sc_hd__a31o_1 _3707_ (.A1(_2856_),
    .A2(_2445_),
    .A3(_2444_),
    .B1(_2443_),
    .X(_2867_));
 sky130_fd_sc_hd__xor2_1 _3708_ (.A(_2866_),
    .B(_2867_),
    .X(_2868_));
 sky130_fd_sc_hd__xnor2_1 _3709_ (.A(_2454_),
    .B(_2868_),
    .Y(_2869_));
 sky130_fd_sc_hd__xnor2_2 _3710_ (.A(_2861_),
    .B(_2869_),
    .Y(_2870_));
 sky130_fd_sc_hd__xnor2_2 _3711_ (.A(_2855_),
    .B(_2870_),
    .Y(_2871_));
 sky130_fd_sc_hd__xnor2_2 _3712_ (.A(_2854_),
    .B(_2871_),
    .Y(_2872_));
 sky130_fd_sc_hd__xor2_2 _3713_ (.A(_2841_),
    .B(_2872_),
    .X(_2873_));
 sky130_fd_sc_hd__xnor2_2 _3714_ (.A(_2839_),
    .B(_2873_),
    .Y(_2874_));
 sky130_fd_sc_hd__xnor2_1 _3715_ (.A(_2832_),
    .B(_2874_),
    .Y(_2875_));
 sky130_fd_sc_hd__xnor2_2 _3716_ (.A(_2830_),
    .B(_2875_),
    .Y(_2876_));
 sky130_fd_sc_hd__xor2_2 _3717_ (.A(_2829_),
    .B(_2876_),
    .X(_2877_));
 sky130_fd_sc_hd__and2_1 _3718_ (.A(net15),
    .B(net14),
    .X(_2878_));
 sky130_fd_sc_hd__clkbuf_4 _3719_ (.A(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__o21ai_1 _3720_ (.A1(_2827_),
    .A2(_2877_),
    .B1(_2879_),
    .Y(_2880_));
 sky130_fd_sc_hd__a21oi_1 _3721_ (.A1(_2827_),
    .A2(_2877_),
    .B1(_2880_),
    .Y(_2881_));
 sky130_fd_sc_hd__clkinv_2 _3722_ (.A(net15),
    .Y(_2882_));
 sky130_fd_sc_hd__clkbuf_4 _3723_ (.A(net14),
    .X(_2883_));
 sky130_fd_sc_hd__nor2_2 _3724_ (.A(_2882_),
    .B(_2883_),
    .Y(_2884_));
 sky130_fd_sc_hd__buf_2 _3725_ (.A(_2884_),
    .X(_2885_));
 sky130_fd_sc_hd__clkbuf_8 _3726_ (.A(\B[2][7] ),
    .X(_2886_));
 sky130_fd_sc_hd__clkbuf_4 _3727_ (.A(\B[0][6] ),
    .X(_2887_));
 sky130_fd_sc_hd__clkbuf_4 _3728_ (.A(_2887_),
    .X(_2888_));
 sky130_fd_sc_hd__and4_1 _3729_ (.A(_2888_),
    .B(_0751_),
    .C(\B[2][0] ),
    .D(_0773_),
    .X(_2889_));
 sky130_fd_sc_hd__a22o_1 _3730_ (.A1(\B[0][7] ),
    .A2(\A[2][0] ),
    .B1(_0872_),
    .B2(\B[0][6] ),
    .X(_2890_));
 sky130_fd_sc_hd__nand4_2 _3731_ (.A(\B[0][6] ),
    .B(\B[0][7] ),
    .C(_0762_),
    .D(_0872_),
    .Y(_2891_));
 sky130_fd_sc_hd__nand4_1 _3732_ (.A(_0806_),
    .B(\B[2][0] ),
    .C(_2890_),
    .D(_2891_),
    .Y(_2892_));
 sky130_fd_sc_hd__a22o_1 _3733_ (.A1(\A[3][7] ),
    .A2(\B[2][0] ),
    .B1(_2890_),
    .B2(_2891_),
    .X(_2893_));
 sky130_fd_sc_hd__nand2_1 _3734_ (.A(\B[0][5] ),
    .B(_0817_),
    .Y(_2894_));
 sky130_fd_sc_hd__buf_2 _3735_ (.A(net59),
    .X(_2895_));
 sky130_fd_sc_hd__clkbuf_4 _3736_ (.A(\B[0][4] ),
    .X(_2896_));
 sky130_fd_sc_hd__a22oi_1 _3737_ (.A1(_2895_),
    .A2(_1004_),
    .B1(_2896_),
    .B2(_0993_),
    .Y(_2897_));
 sky130_fd_sc_hd__and4_1 _3738_ (.A(_0960_),
    .B(_2895_),
    .C(_0905_),
    .D(_2896_),
    .X(_2898_));
 sky130_fd_sc_hd__o21bai_1 _3739_ (.A1(_2894_),
    .A2(_2897_),
    .B1_N(_2898_),
    .Y(_2899_));
 sky130_fd_sc_hd__a21o_1 _3740_ (.A1(_2892_),
    .A2(_2893_),
    .B1(_2899_),
    .X(_2900_));
 sky130_fd_sc_hd__nand3_1 _3741_ (.A(_2899_),
    .B(_2892_),
    .C(_2893_),
    .Y(_2901_));
 sky130_fd_sc_hd__a21bo_1 _3742_ (.A1(_2889_),
    .A2(_2900_),
    .B1_N(_2901_),
    .X(_2902_));
 sky130_fd_sc_hd__clkbuf_4 _3743_ (.A(\B[2][1] ),
    .X(_2903_));
 sky130_fd_sc_hd__a22o_1 _3744_ (.A1(\A[3][7] ),
    .A2(_2903_),
    .B1(\B[2][2] ),
    .B2(\A[3][6] ),
    .X(_2904_));
 sky130_fd_sc_hd__clkbuf_4 _3745_ (.A(\B[2][2] ),
    .X(_2905_));
 sky130_fd_sc_hd__nand4_1 _3746_ (.A(\A[3][7] ),
    .B(_1114_),
    .C(_2903_),
    .D(_2905_),
    .Y(_2906_));
 sky130_fd_sc_hd__and2_1 _3747_ (.A(_1158_),
    .B(\B[2][3] ),
    .X(_2907_));
 sky130_fd_sc_hd__nand3_1 _3748_ (.A(_2904_),
    .B(_2906_),
    .C(_2907_),
    .Y(_2908_));
 sky130_fd_sc_hd__a21o_1 _3749_ (.A1(_2904_),
    .A2(_2906_),
    .B1(_2907_),
    .X(_2909_));
 sky130_fd_sc_hd__nand2_1 _3750_ (.A(\B[2][3] ),
    .B(_1466_),
    .Y(_2910_));
 sky130_fd_sc_hd__a22oi_2 _3751_ (.A1(_1114_),
    .A2(_2903_),
    .B1(_2905_),
    .B2(_1158_),
    .Y(_2911_));
 sky130_fd_sc_hd__and4_1 _3752_ (.A(\A[3][6] ),
    .B(\A[3][5] ),
    .C(\B[2][1] ),
    .D(\B[2][2] ),
    .X(_2912_));
 sky130_fd_sc_hd__o21bai_1 _3753_ (.A1(_2910_),
    .A2(_2911_),
    .B1_N(_2912_),
    .Y(_2913_));
 sky130_fd_sc_hd__and3_1 _3754_ (.A(_2908_),
    .B(_2909_),
    .C(_2913_),
    .X(_2914_));
 sky130_fd_sc_hd__a21oi_1 _3755_ (.A1(_2908_),
    .A2(_2909_),
    .B1(_2913_),
    .Y(_2915_));
 sky130_fd_sc_hd__clkbuf_4 _3756_ (.A(\B[2][5] ),
    .X(_2916_));
 sky130_fd_sc_hd__buf_4 _3757_ (.A(\B[2][4] ),
    .X(_2917_));
 sky130_fd_sc_hd__a22oi_1 _3758_ (.A1(_2916_),
    .A2(_1323_),
    .B1(_2917_),
    .B2(_1213_),
    .Y(_2918_));
 sky130_fd_sc_hd__and4_1 _3759_ (.A(\B[2][5] ),
    .B(\A[3][3] ),
    .C(\B[2][4] ),
    .D(_1466_),
    .X(_2919_));
 sky130_fd_sc_hd__nor2_1 _3760_ (.A(_2918_),
    .B(_2919_),
    .Y(_2920_));
 sky130_fd_sc_hd__buf_4 _3761_ (.A(net48),
    .X(_2921_));
 sky130_fd_sc_hd__nand2_1 _3762_ (.A(_2921_),
    .B(_0707_),
    .Y(_2922_));
 sky130_fd_sc_hd__xnor2_1 _3763_ (.A(_2920_),
    .B(_2922_),
    .Y(_2923_));
 sky130_fd_sc_hd__or3b_1 _3764_ (.A(_2914_),
    .B(_2915_),
    .C_N(_2923_),
    .X(_2924_));
 sky130_fd_sc_hd__o21bai_1 _3765_ (.A1(_2914_),
    .A2(_2915_),
    .B1_N(_2923_),
    .Y(_2925_));
 sky130_fd_sc_hd__and3_1 _3766_ (.A(_2902_),
    .B(_2924_),
    .C(_2925_),
    .X(_2926_));
 sky130_fd_sc_hd__or3_1 _3767_ (.A(_2912_),
    .B(_2910_),
    .C(_2911_),
    .X(_2927_));
 sky130_fd_sc_hd__o21ai_1 _3768_ (.A1(_2912_),
    .A2(_2911_),
    .B1(_2910_),
    .Y(_2928_));
 sky130_fd_sc_hd__nand2_1 _3769_ (.A(\B[2][3] ),
    .B(_1323_),
    .Y(_2929_));
 sky130_fd_sc_hd__a22oi_2 _3770_ (.A1(_1158_),
    .A2(_2903_),
    .B1(_2905_),
    .B2(_1466_),
    .Y(_2930_));
 sky130_fd_sc_hd__and4_1 _3771_ (.A(_1158_),
    .B(\B[2][1] ),
    .C(\B[2][2] ),
    .D(_1466_),
    .X(_2931_));
 sky130_fd_sc_hd__o21bai_1 _3772_ (.A1(_2929_),
    .A2(_2930_),
    .B1_N(_2931_),
    .Y(_2932_));
 sky130_fd_sc_hd__nand3_2 _3773_ (.A(_2927_),
    .B(_2928_),
    .C(_2932_),
    .Y(_2933_));
 sky130_fd_sc_hd__a22oi_1 _3774_ (.A1(_2916_),
    .A2(_0707_),
    .B1(_1323_),
    .B2(_2917_),
    .Y(_2934_));
 sky130_fd_sc_hd__and4_1 _3775_ (.A(_2916_),
    .B(_2559_),
    .C(_1323_),
    .D(\B[2][4] ),
    .X(_2935_));
 sky130_fd_sc_hd__nor2_1 _3776_ (.A(_2934_),
    .B(_2935_),
    .Y(_2936_));
 sky130_fd_sc_hd__nand2_1 _3777_ (.A(_2921_),
    .B(_1609_),
    .Y(_2937_));
 sky130_fd_sc_hd__xnor2_1 _3778_ (.A(_2936_),
    .B(_2937_),
    .Y(_2938_));
 sky130_fd_sc_hd__a21o_1 _3779_ (.A1(_2927_),
    .A2(_2928_),
    .B1(_2932_),
    .X(_2939_));
 sky130_fd_sc_hd__nand3_1 _3780_ (.A(_2933_),
    .B(_2938_),
    .C(_2939_),
    .Y(_2940_));
 sky130_fd_sc_hd__a21oi_1 _3781_ (.A1(_2924_),
    .A2(_2925_),
    .B1(_2902_),
    .Y(_2941_));
 sky130_fd_sc_hd__a211oi_1 _3782_ (.A1(_2933_),
    .A2(_2940_),
    .B1(_2941_),
    .C1(_2926_),
    .Y(_2942_));
 sky130_fd_sc_hd__o21ba_1 _3783_ (.A1(_2918_),
    .A2(_2922_),
    .B1_N(_2919_),
    .X(_2943_));
 sky130_fd_sc_hd__o21ba_1 _3784_ (.A1(_2926_),
    .A2(_2942_),
    .B1_N(_2943_),
    .X(_2944_));
 sky130_fd_sc_hd__or3b_1 _3785_ (.A(_2926_),
    .B(_2942_),
    .C_N(_2943_),
    .X(_2945_));
 sky130_fd_sc_hd__and2b_1 _3786_ (.A_N(_2944_),
    .B(_2945_),
    .X(_2946_));
 sky130_fd_sc_hd__a31o_2 _3787_ (.A1(_2886_),
    .A2(_0718_),
    .A3(_2946_),
    .B1(_2944_),
    .X(_2947_));
 sky130_fd_sc_hd__a22oi_1 _3788_ (.A1(_1740_),
    .A2(\B[2][4] ),
    .B1(_1213_),
    .B2(_2916_),
    .Y(_2948_));
 sky130_fd_sc_hd__and4_1 _3789_ (.A(\B[2][5] ),
    .B(_1158_),
    .C(\B[2][4] ),
    .D(_1466_),
    .X(_2949_));
 sky130_fd_sc_hd__nor2_1 _3790_ (.A(_2948_),
    .B(_2949_),
    .Y(_2950_));
 sky130_fd_sc_hd__nand2_1 _3791_ (.A(_2921_),
    .B(_1532_),
    .Y(_2951_));
 sky130_fd_sc_hd__xnor2_1 _3792_ (.A(_2950_),
    .B(_2951_),
    .Y(_2952_));
 sky130_fd_sc_hd__nand2_1 _3793_ (.A(_1114_),
    .B(_2905_),
    .Y(_2953_));
 sky130_fd_sc_hd__nand2_1 _3794_ (.A(\A[3][7] ),
    .B(\B[2][3] ),
    .Y(_2954_));
 sky130_fd_sc_hd__a22o_1 _3795_ (.A1(\A[3][7] ),
    .A2(_2905_),
    .B1(\B[2][3] ),
    .B2(_1114_),
    .X(_2955_));
 sky130_fd_sc_hd__o21a_1 _3796_ (.A1(_2953_),
    .A2(_2954_),
    .B1(_2955_),
    .X(_2956_));
 sky130_fd_sc_hd__a21boi_2 _3797_ (.A1(_2904_),
    .A2(_2907_),
    .B1_N(_2906_),
    .Y(_2957_));
 sky130_fd_sc_hd__xnor2_1 _3798_ (.A(_2956_),
    .B(_2957_),
    .Y(_2958_));
 sky130_fd_sc_hd__xnor2_1 _3799_ (.A(_2952_),
    .B(_2958_),
    .Y(_2959_));
 sky130_fd_sc_hd__nand2_1 _3800_ (.A(_2891_),
    .B(_2892_),
    .Y(_2960_));
 sky130_fd_sc_hd__a22o_1 _3801_ (.A1(_0905_),
    .A2(_2896_),
    .B1(_2238_),
    .B2(_2895_),
    .X(_2961_));
 sky130_fd_sc_hd__and4_1 _3802_ (.A(_2895_),
    .B(_0905_),
    .C(\B[0][4] ),
    .D(_2238_),
    .X(_2962_));
 sky130_fd_sc_hd__a31oi_2 _3803_ (.A1(\B[0][5] ),
    .A2(_0971_),
    .A3(_2961_),
    .B1(_2962_),
    .Y(_2963_));
 sky130_fd_sc_hd__clkbuf_4 _3804_ (.A(\B[0][7] ),
    .X(_2964_));
 sky130_fd_sc_hd__a22oi_2 _3805_ (.A1(_2964_),
    .A2(_0817_),
    .B1(_0971_),
    .B2(_2887_),
    .Y(_2965_));
 sky130_fd_sc_hd__and4_1 _3806_ (.A(\B[0][6] ),
    .B(\B[0][7] ),
    .C(_0817_),
    .D(_0993_),
    .X(_2966_));
 sky130_fd_sc_hd__nor2_1 _3807_ (.A(_2965_),
    .B(_2966_),
    .Y(_2967_));
 sky130_fd_sc_hd__xnor2_2 _3808_ (.A(_2963_),
    .B(_2967_),
    .Y(_2968_));
 sky130_fd_sc_hd__or3_1 _3809_ (.A(_2963_),
    .B(_2965_),
    .C(_2966_),
    .X(_2969_));
 sky130_fd_sc_hd__a21bo_1 _3810_ (.A1(_2960_),
    .A2(_2968_),
    .B1_N(_2969_),
    .X(_2970_));
 sky130_fd_sc_hd__and2b_1 _3811_ (.A_N(_2959_),
    .B(_2970_),
    .X(_2971_));
 sky130_fd_sc_hd__nor3b_1 _3812_ (.A(_2914_),
    .B(_2915_),
    .C_N(_2923_),
    .Y(_2972_));
 sky130_fd_sc_hd__xnor2_1 _3813_ (.A(_2970_),
    .B(_2959_),
    .Y(_2973_));
 sky130_fd_sc_hd__o21a_1 _3814_ (.A1(_2914_),
    .A2(_2972_),
    .B1(_2973_),
    .X(_2974_));
 sky130_fd_sc_hd__o21ba_1 _3815_ (.A1(_2948_),
    .A2(_2951_),
    .B1_N(_2949_),
    .X(_2975_));
 sky130_fd_sc_hd__o21ba_1 _3816_ (.A1(_2971_),
    .A2(_2974_),
    .B1_N(_2975_),
    .X(_2976_));
 sky130_fd_sc_hd__or3b_1 _3817_ (.A(_2971_),
    .B(_2974_),
    .C_N(_2975_),
    .X(_2977_));
 sky130_fd_sc_hd__and2b_2 _3818_ (.A_N(_2976_),
    .B(_2977_),
    .X(_2978_));
 sky130_fd_sc_hd__nand2_1 _3819_ (.A(\B[2][7] ),
    .B(_1532_),
    .Y(_2979_));
 sky130_fd_sc_hd__xnor2_4 _3820_ (.A(_2978_),
    .B(_2979_),
    .Y(_2980_));
 sky130_fd_sc_hd__inv_2 _3821_ (.A(_2955_),
    .Y(_2981_));
 sky130_fd_sc_hd__nor2_1 _3822_ (.A(_2953_),
    .B(_2954_),
    .Y(_2982_));
 sky130_fd_sc_hd__nand2_1 _3823_ (.A(_2952_),
    .B(_2958_),
    .Y(_2983_));
 sky130_fd_sc_hd__o31ai_4 _3824_ (.A1(_2981_),
    .A2(_2982_),
    .A3(_2957_),
    .B1(_2983_),
    .Y(_2984_));
 sky130_fd_sc_hd__a22oi_1 _3825_ (.A1(\B[0][7] ),
    .A2(_0993_),
    .B1(_0916_),
    .B2(_2887_),
    .Y(_2985_));
 sky130_fd_sc_hd__and4_1 _3826_ (.A(\B[0][6] ),
    .B(\B[0][7] ),
    .C(_0993_),
    .D(_1004_),
    .X(_2986_));
 sky130_fd_sc_hd__or2_1 _3827_ (.A(_2985_),
    .B(_2986_),
    .X(_2987_));
 sky130_fd_sc_hd__buf_4 _3828_ (.A(\B[0][5] ),
    .X(_2988_));
 sky130_fd_sc_hd__a22o_1 _3829_ (.A1(_2526_),
    .A2(\B[0][3] ),
    .B1(_2896_),
    .B2(\A[2][4] ),
    .X(_2989_));
 sky130_fd_sc_hd__and4_1 _3830_ (.A(_2526_),
    .B(\B[0][3] ),
    .C(\B[0][4] ),
    .D(\A[2][4] ),
    .X(_2990_));
 sky130_fd_sc_hd__a31o_1 _3831_ (.A1(_2988_),
    .A2(_0916_),
    .A3(_2989_),
    .B1(_2990_),
    .X(_2991_));
 sky130_fd_sc_hd__or2b_1 _3832_ (.A(_2987_),
    .B_N(_2991_),
    .X(_2992_));
 sky130_fd_sc_hd__xnor2_1 _3833_ (.A(_2991_),
    .B(_2987_),
    .Y(_2993_));
 sky130_fd_sc_hd__nand2_1 _3834_ (.A(_2966_),
    .B(_2993_),
    .Y(_2994_));
 sky130_fd_sc_hd__a22o_1 _3835_ (.A1(_2916_),
    .A2(_1740_),
    .B1(_2917_),
    .B2(_1114_),
    .X(_2995_));
 sky130_fd_sc_hd__nand4_1 _3836_ (.A(_2916_),
    .B(_0751_),
    .C(_1740_),
    .D(_2917_),
    .Y(_2996_));
 sky130_fd_sc_hd__and2_1 _3837_ (.A(\B[2][6] ),
    .B(_1213_),
    .X(_2997_));
 sky130_fd_sc_hd__a21oi_1 _3838_ (.A1(_2995_),
    .A2(_2996_),
    .B1(_2997_),
    .Y(_2998_));
 sky130_fd_sc_hd__and3_1 _3839_ (.A(_2995_),
    .B(_2996_),
    .C(_2997_),
    .X(_2999_));
 sky130_fd_sc_hd__nor2_1 _3840_ (.A(_2998_),
    .B(_2999_),
    .Y(_3000_));
 sky130_fd_sc_hd__clkbuf_4 _3841_ (.A(\B[2][3] ),
    .X(_3001_));
 sky130_fd_sc_hd__buf_4 _3842_ (.A(_3001_),
    .X(_3002_));
 sky130_fd_sc_hd__and3_1 _3843_ (.A(_0806_),
    .B(_3002_),
    .C(_2953_),
    .X(_3003_));
 sky130_fd_sc_hd__xnor2_2 _3844_ (.A(_3000_),
    .B(_3003_),
    .Y(_3004_));
 sky130_fd_sc_hd__a21oi_1 _3845_ (.A1(_2992_),
    .A2(_2994_),
    .B1(_3004_),
    .Y(_3005_));
 sky130_fd_sc_hd__nand3_1 _3846_ (.A(_2992_),
    .B(_2994_),
    .C(_3004_),
    .Y(_3006_));
 sky130_fd_sc_hd__and2b_1 _3847_ (.A_N(_3005_),
    .B(_3006_),
    .X(_3007_));
 sky130_fd_sc_hd__xor2_4 _3848_ (.A(_2984_),
    .B(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__a22o_1 _3849_ (.A1(\A[2][6] ),
    .A2(\B[0][3] ),
    .B1(\B[0][4] ),
    .B2(_2526_),
    .X(_3009_));
 sky130_fd_sc_hd__nand4_1 _3850_ (.A(_2392_),
    .B(_2526_),
    .C(_2895_),
    .D(_2896_),
    .Y(_3010_));
 sky130_fd_sc_hd__and2_1 _3851_ (.A(\B[0][5] ),
    .B(\A[2][4] ),
    .X(_3011_));
 sky130_fd_sc_hd__a21o_1 _3852_ (.A1(_3009_),
    .A2(_3010_),
    .B1(_3011_),
    .X(_3012_));
 sky130_fd_sc_hd__nand3_1 _3853_ (.A(_3009_),
    .B(_3010_),
    .C(_3011_),
    .Y(_3013_));
 sky130_fd_sc_hd__clkbuf_4 _3854_ (.A(net54),
    .X(_3014_));
 sky130_fd_sc_hd__clkbuf_4 _3855_ (.A(\B[0][1] ),
    .X(_3015_));
 sky130_fd_sc_hd__nand2_1 _3856_ (.A(_2392_),
    .B(_3015_),
    .Y(_3016_));
 sky130_fd_sc_hd__and3_1 _3857_ (.A(_2431_),
    .B(_3014_),
    .C(_3016_),
    .X(_3017_));
 sky130_fd_sc_hd__and3_1 _3858_ (.A(_3012_),
    .B(_3013_),
    .C(_3017_),
    .X(_3018_));
 sky130_fd_sc_hd__and4_1 _3859_ (.A(\A[2][7] ),
    .B(\A[2][6] ),
    .C(\B[0][1] ),
    .D(\B[0][2] ),
    .X(_3019_));
 sky130_fd_sc_hd__nand2_1 _3860_ (.A(_2431_),
    .B(_2895_),
    .Y(_3020_));
 sky130_fd_sc_hd__nand2_1 _3861_ (.A(_2392_),
    .B(_2896_),
    .Y(_3021_));
 sky130_fd_sc_hd__and4_1 _3862_ (.A(\A[2][7] ),
    .B(\A[2][6] ),
    .C(_2895_),
    .D(_2896_),
    .X(_3022_));
 sky130_fd_sc_hd__a21oi_1 _3863_ (.A1(_3020_),
    .A2(_3021_),
    .B1(_3022_),
    .Y(_3023_));
 sky130_fd_sc_hd__nand2_1 _3864_ (.A(_2988_),
    .B(_2218_),
    .Y(_3024_));
 sky130_fd_sc_hd__xnor2_1 _3865_ (.A(_3023_),
    .B(_3024_),
    .Y(_3025_));
 sky130_fd_sc_hd__o21a_1 _3866_ (.A1(_3018_),
    .A2(_3019_),
    .B1(_3025_),
    .X(_3026_));
 sky130_fd_sc_hd__or3_1 _3867_ (.A(_3025_),
    .B(_3018_),
    .C(_3019_),
    .X(_3027_));
 sky130_fd_sc_hd__and2b_1 _3868_ (.A_N(_3026_),
    .B(_3027_),
    .X(_3028_));
 sky130_fd_sc_hd__a21bo_1 _3869_ (.A1(_3009_),
    .A2(_3011_),
    .B1_N(_3010_),
    .X(_3029_));
 sky130_fd_sc_hd__nand2_1 _3870_ (.A(_2964_),
    .B(_0916_),
    .Y(_3030_));
 sky130_fd_sc_hd__nand2_1 _3871_ (.A(_2887_),
    .B(_1915_),
    .Y(_3031_));
 sky130_fd_sc_hd__and4_1 _3872_ (.A(\B[0][6] ),
    .B(\B[0][7] ),
    .C(_1004_),
    .D(_2238_),
    .X(_3032_));
 sky130_fd_sc_hd__a21o_1 _3873_ (.A1(_3030_),
    .A2(_3031_),
    .B1(_3032_),
    .X(_3033_));
 sky130_fd_sc_hd__xnor2_1 _3874_ (.A(_3029_),
    .B(_3033_),
    .Y(_3034_));
 sky130_fd_sc_hd__nor2_1 _3875_ (.A(_2986_),
    .B(_3034_),
    .Y(_3035_));
 sky130_fd_sc_hd__and2_1 _3876_ (.A(_2986_),
    .B(_3034_),
    .X(_3036_));
 sky130_fd_sc_hd__nor2_2 _3877_ (.A(_3035_),
    .B(_3036_),
    .Y(_3037_));
 sky130_fd_sc_hd__xor2_4 _3878_ (.A(_3028_),
    .B(_3037_),
    .X(_3038_));
 sky130_fd_sc_hd__a21oi_2 _3879_ (.A1(_3012_),
    .A2(_3013_),
    .B1(_3017_),
    .Y(_3039_));
 sky130_fd_sc_hd__and2b_1 _3880_ (.A_N(_2990_),
    .B(_2989_),
    .X(_3040_));
 sky130_fd_sc_hd__nand2_1 _3881_ (.A(_2988_),
    .B(_0916_),
    .Y(_3041_));
 sky130_fd_sc_hd__xnor2_2 _3882_ (.A(_3040_),
    .B(_3041_),
    .Y(_3042_));
 sky130_fd_sc_hd__a22oi_1 _3883_ (.A1(\A[2][7] ),
    .A2(_3015_),
    .B1(_3014_),
    .B2(_2392_),
    .Y(_3043_));
 sky130_fd_sc_hd__or2_1 _3884_ (.A(_3019_),
    .B(_3043_),
    .X(_3044_));
 sky130_fd_sc_hd__and2_1 _3885_ (.A(_2526_),
    .B(\B[0][2] ),
    .X(_3045_));
 sky130_fd_sc_hd__clkbuf_4 _3886_ (.A(\B[0][0] ),
    .X(_3046_));
 sky130_fd_sc_hd__a22o_1 _3887_ (.A1(\A[2][7] ),
    .A2(_3046_),
    .B1(_3015_),
    .B2(_2392_),
    .X(_3047_));
 sky130_fd_sc_hd__nand4_1 _3888_ (.A(\A[2][7] ),
    .B(_2392_),
    .C(_3046_),
    .D(_3015_),
    .Y(_3048_));
 sky130_fd_sc_hd__a21bo_1 _3889_ (.A1(_3045_),
    .A2(_3047_),
    .B1_N(_3048_),
    .X(_3049_));
 sky130_fd_sc_hd__xnor2_2 _3890_ (.A(_3044_),
    .B(_3049_),
    .Y(_3050_));
 sky130_fd_sc_hd__or2b_1 _3891_ (.A(_3044_),
    .B_N(_3049_),
    .X(_3051_));
 sky130_fd_sc_hd__a21boi_4 _3892_ (.A1(_3042_),
    .A2(_3050_),
    .B1_N(_3051_),
    .Y(_3052_));
 sky130_fd_sc_hd__or2_1 _3893_ (.A(_2966_),
    .B(_2993_),
    .X(_3053_));
 sky130_fd_sc_hd__nand2_2 _3894_ (.A(_2994_),
    .B(_3053_),
    .Y(_3054_));
 sky130_fd_sc_hd__or2_2 _3895_ (.A(_3018_),
    .B(_3039_),
    .X(_3055_));
 sky130_fd_sc_hd__xnor2_4 _3896_ (.A(_3055_),
    .B(_3052_),
    .Y(_3056_));
 sky130_fd_sc_hd__o32ai_4 _3897_ (.A1(_3018_),
    .A2(_3039_),
    .A3(_3052_),
    .B1(_3054_),
    .B2(_3056_),
    .Y(_3057_));
 sky130_fd_sc_hd__xor2_4 _3898_ (.A(_3038_),
    .B(_3057_),
    .X(_3058_));
 sky130_fd_sc_hd__xnor2_4 _3899_ (.A(_3008_),
    .B(_3058_),
    .Y(_3059_));
 sky130_fd_sc_hd__nor3_1 _3900_ (.A(_2914_),
    .B(_2972_),
    .C(_2973_),
    .Y(_3060_));
 sky130_fd_sc_hd__nor2_1 _3901_ (.A(_2974_),
    .B(_3060_),
    .Y(_3061_));
 sky130_fd_sc_hd__xor2_4 _3902_ (.A(_3054_),
    .B(_3056_),
    .X(_3062_));
 sky130_fd_sc_hd__xnor2_2 _3903_ (.A(_2960_),
    .B(_2968_),
    .Y(_3063_));
 sky130_fd_sc_hd__xnor2_2 _3904_ (.A(_3042_),
    .B(_3050_),
    .Y(_3064_));
 sky130_fd_sc_hd__nand2_1 _3905_ (.A(_2988_),
    .B(_0971_),
    .Y(_3065_));
 sky130_fd_sc_hd__and2b_1 _3906_ (.A_N(_2962_),
    .B(_2961_),
    .X(_3066_));
 sky130_fd_sc_hd__xnor2_1 _3907_ (.A(_3065_),
    .B(_3066_),
    .Y(_3067_));
 sky130_fd_sc_hd__nand3_1 _3908_ (.A(_3048_),
    .B(_3045_),
    .C(_3047_),
    .Y(_3068_));
 sky130_fd_sc_hd__a21o_1 _3909_ (.A1(_3048_),
    .A2(_3047_),
    .B1(_3045_),
    .X(_3069_));
 sky130_fd_sc_hd__nand2_1 _3910_ (.A(_3014_),
    .B(_2238_),
    .Y(_3070_));
 sky130_fd_sc_hd__a22oi_2 _3911_ (.A1(_2392_),
    .A2(_3046_),
    .B1(_3015_),
    .B2(_2526_),
    .Y(_3071_));
 sky130_fd_sc_hd__and4_1 _3912_ (.A(\A[2][6] ),
    .B(_2526_),
    .C(\B[0][0] ),
    .D(\B[0][1] ),
    .X(_3072_));
 sky130_fd_sc_hd__o21bai_1 _3913_ (.A1(_3070_),
    .A2(_3071_),
    .B1_N(_3072_),
    .Y(_3073_));
 sky130_fd_sc_hd__a21o_1 _3914_ (.A1(_3068_),
    .A2(_3069_),
    .B1(_3073_),
    .X(_3074_));
 sky130_fd_sc_hd__nand3_1 _3915_ (.A(_3068_),
    .B(_3069_),
    .C(_3073_),
    .Y(_3075_));
 sky130_fd_sc_hd__a21bo_1 _3916_ (.A1(_3067_),
    .A2(_3074_),
    .B1_N(_3075_),
    .X(_3076_));
 sky130_fd_sc_hd__xor2_2 _3917_ (.A(_3064_),
    .B(_3076_),
    .X(_3077_));
 sky130_fd_sc_hd__or2b_1 _3918_ (.A(_3064_),
    .B_N(_3076_),
    .X(_3078_));
 sky130_fd_sc_hd__o21a_1 _3919_ (.A1(_3063_),
    .A2(_3077_),
    .B1(_3078_),
    .X(_3079_));
 sky130_fd_sc_hd__xnor2_4 _3920_ (.A(_3062_),
    .B(_3079_),
    .Y(_3080_));
 sky130_fd_sc_hd__or2b_1 _3921_ (.A(_3079_),
    .B_N(_3062_),
    .X(_3081_));
 sky130_fd_sc_hd__a21boi_2 _3922_ (.A1(_3061_),
    .A2(_3080_),
    .B1_N(_3081_),
    .Y(_3082_));
 sky130_fd_sc_hd__xor2_4 _3923_ (.A(_3059_),
    .B(_3082_),
    .X(_3083_));
 sky130_fd_sc_hd__xnor2_4 _3924_ (.A(_2980_),
    .B(_3083_),
    .Y(_3084_));
 sky130_fd_sc_hd__nand2_1 _3925_ (.A(\B[2][7] ),
    .B(_0718_),
    .Y(_3085_));
 sky130_fd_sc_hd__xnor2_2 _3926_ (.A(_2946_),
    .B(_3085_),
    .Y(_3086_));
 sky130_fd_sc_hd__xnor2_2 _3927_ (.A(_3061_),
    .B(_3080_),
    .Y(_3087_));
 sky130_fd_sc_hd__o211a_1 _3928_ (.A1(_2926_),
    .A2(_2941_),
    .B1(_2940_),
    .C1(_2933_),
    .X(_3088_));
 sky130_fd_sc_hd__nor2_1 _3929_ (.A(_2942_),
    .B(_3088_),
    .Y(_3089_));
 sky130_fd_sc_hd__xnor2_2 _3930_ (.A(_3063_),
    .B(_3077_),
    .Y(_3090_));
 sky130_fd_sc_hd__and3_1 _3931_ (.A(_2901_),
    .B(_2889_),
    .C(_2900_),
    .X(_3091_));
 sky130_fd_sc_hd__a21oi_1 _3932_ (.A1(_2901_),
    .A2(_2900_),
    .B1(_2889_),
    .Y(_3092_));
 sky130_fd_sc_hd__or2_1 _3933_ (.A(_3091_),
    .B(_3092_),
    .X(_3093_));
 sky130_fd_sc_hd__nand3_1 _3934_ (.A(_3075_),
    .B(_3067_),
    .C(_3074_),
    .Y(_3094_));
 sky130_fd_sc_hd__a21o_1 _3935_ (.A1(_3075_),
    .A2(_3074_),
    .B1(_3067_),
    .X(_3095_));
 sky130_fd_sc_hd__nor2_1 _3936_ (.A(_2898_),
    .B(_2897_),
    .Y(_3096_));
 sky130_fd_sc_hd__xnor2_1 _3937_ (.A(_2894_),
    .B(_3096_),
    .Y(_3097_));
 sky130_fd_sc_hd__or3_1 _3938_ (.A(_3072_),
    .B(_3070_),
    .C(_3071_),
    .X(_3098_));
 sky130_fd_sc_hd__o21ai_1 _3939_ (.A1(_3072_),
    .A2(_3071_),
    .B1(_3070_),
    .Y(_3099_));
 sky130_fd_sc_hd__nand2_1 _3940_ (.A(_3014_),
    .B(_0905_),
    .Y(_3100_));
 sky130_fd_sc_hd__a22oi_2 _3941_ (.A1(_2526_),
    .A2(\B[0][0] ),
    .B1(_3015_),
    .B2(_2238_),
    .Y(_3101_));
 sky130_fd_sc_hd__and4_1 _3942_ (.A(_2526_),
    .B(\B[0][0] ),
    .C(\B[0][1] ),
    .D(\A[2][4] ),
    .X(_3102_));
 sky130_fd_sc_hd__o21bai_1 _3943_ (.A1(_3100_),
    .A2(_3101_),
    .B1_N(_3102_),
    .Y(_0064_));
 sky130_fd_sc_hd__a21o_1 _3944_ (.A1(_3098_),
    .A2(_3099_),
    .B1(_0064_),
    .X(_0065_));
 sky130_fd_sc_hd__nand3_1 _3945_ (.A(_3098_),
    .B(_3099_),
    .C(_0064_),
    .Y(_0066_));
 sky130_fd_sc_hd__a21bo_1 _3946_ (.A1(_3097_),
    .A2(_0065_),
    .B1_N(_0066_),
    .X(_0067_));
 sky130_fd_sc_hd__a21oi_1 _3947_ (.A1(_3094_),
    .A2(_3095_),
    .B1(_0067_),
    .Y(_0068_));
 sky130_fd_sc_hd__and3_1 _3948_ (.A(_3094_),
    .B(_3095_),
    .C(_0067_),
    .X(_0069_));
 sky130_fd_sc_hd__o21ba_1 _3949_ (.A1(_3093_),
    .A2(_0068_),
    .B1_N(_0069_),
    .X(_0070_));
 sky130_fd_sc_hd__xor2_2 _3950_ (.A(_3090_),
    .B(_0070_),
    .X(_0071_));
 sky130_fd_sc_hd__nor2_1 _3951_ (.A(_3090_),
    .B(_0070_),
    .Y(_0072_));
 sky130_fd_sc_hd__a21o_1 _3952_ (.A1(_3089_),
    .A2(_0071_),
    .B1(_0072_),
    .X(_0073_));
 sky130_fd_sc_hd__xnor2_2 _3953_ (.A(_3087_),
    .B(_0073_),
    .Y(_0074_));
 sky130_fd_sc_hd__or2b_1 _3954_ (.A(_3087_),
    .B_N(_0073_),
    .X(_0075_));
 sky130_fd_sc_hd__a21boi_2 _3955_ (.A1(_3086_),
    .A2(_0074_),
    .B1_N(_0075_),
    .Y(_0076_));
 sky130_fd_sc_hd__xor2_4 _3956_ (.A(_3084_),
    .B(_0076_),
    .X(_0077_));
 sky130_fd_sc_hd__xnor2_4 _3957_ (.A(_2947_),
    .B(_0077_),
    .Y(_0078_));
 sky130_fd_sc_hd__buf_4 _3958_ (.A(_2886_),
    .X(_0079_));
 sky130_fd_sc_hd__and4_1 _3959_ (.A(_0872_),
    .B(\A[2][2] ),
    .C(\B[0][3] ),
    .D(\B[0][4] ),
    .X(_0080_));
 sky130_fd_sc_hd__nand2_1 _3960_ (.A(\B[0][5] ),
    .B(_0762_),
    .Y(_0081_));
 sky130_fd_sc_hd__a22oi_1 _3961_ (.A1(_0993_),
    .A2(_2895_),
    .B1(_2896_),
    .B2(_0817_),
    .Y(_0082_));
 sky130_fd_sc_hd__or2_1 _3962_ (.A(_0082_),
    .B(_0080_),
    .X(_0083_));
 sky130_fd_sc_hd__nor2_1 _3963_ (.A(_0081_),
    .B(_0083_),
    .Y(_0084_));
 sky130_fd_sc_hd__buf_4 _3964_ (.A(\B[2][0] ),
    .X(_0085_));
 sky130_fd_sc_hd__a22oi_1 _3965_ (.A1(_0751_),
    .A2(_0085_),
    .B1(_0773_),
    .B2(_2888_),
    .Y(_0086_));
 sky130_fd_sc_hd__nor2_1 _3966_ (.A(_2889_),
    .B(_0086_),
    .Y(_0087_));
 sky130_fd_sc_hd__o21a_2 _3967_ (.A1(_0080_),
    .A2(_0084_),
    .B1(_0087_),
    .X(_0088_));
 sky130_fd_sc_hd__a21o_1 _3968_ (.A1(_2933_),
    .A2(_2939_),
    .B1(_2938_),
    .X(_0089_));
 sky130_fd_sc_hd__and3_1 _3969_ (.A(_2940_),
    .B(_0088_),
    .C(_0089_),
    .X(_0090_));
 sky130_fd_sc_hd__or3_1 _3970_ (.A(_2931_),
    .B(_2929_),
    .C(_2930_),
    .X(_0091_));
 sky130_fd_sc_hd__o21ai_1 _3971_ (.A1(_2931_),
    .A2(_2930_),
    .B1(_2929_),
    .Y(_0092_));
 sky130_fd_sc_hd__nand2_1 _3972_ (.A(_2559_),
    .B(\B[2][3] ),
    .Y(_0093_));
 sky130_fd_sc_hd__a22oi_2 _3973_ (.A1(\B[2][2] ),
    .A2(\A[3][3] ),
    .B1(_1466_),
    .B2(_2903_),
    .Y(_0094_));
 sky130_fd_sc_hd__and4_1 _3974_ (.A(\B[2][1] ),
    .B(\B[2][2] ),
    .C(\A[3][3] ),
    .D(\A[3][4] ),
    .X(_0095_));
 sky130_fd_sc_hd__o21bai_1 _3975_ (.A1(_0093_),
    .A2(_0094_),
    .B1_N(_0095_),
    .Y(_0096_));
 sky130_fd_sc_hd__nand3_1 _3976_ (.A(_0091_),
    .B(_0092_),
    .C(_0096_),
    .Y(_0097_));
 sky130_fd_sc_hd__a22oi_1 _3977_ (.A1(_2916_),
    .A2(_1598_),
    .B1(_0707_),
    .B2(_2917_),
    .Y(_0098_));
 sky130_fd_sc_hd__and4_1 _3978_ (.A(_2916_),
    .B(\A[3][1] ),
    .C(_2559_),
    .D(\B[2][4] ),
    .X(_0099_));
 sky130_fd_sc_hd__nor2_1 _3979_ (.A(_0098_),
    .B(_0099_),
    .Y(_0100_));
 sky130_fd_sc_hd__nand2_1 _3980_ (.A(_2921_),
    .B(_2568_),
    .Y(_0101_));
 sky130_fd_sc_hd__xnor2_1 _3981_ (.A(_0100_),
    .B(_0101_),
    .Y(_0102_));
 sky130_fd_sc_hd__a21o_1 _3982_ (.A1(_0091_),
    .A2(_0092_),
    .B1(_0096_),
    .X(_0103_));
 sky130_fd_sc_hd__nand3_1 _3983_ (.A(_0097_),
    .B(_0102_),
    .C(_0103_),
    .Y(_0104_));
 sky130_fd_sc_hd__nand2_1 _3984_ (.A(_0097_),
    .B(_0104_),
    .Y(_0105_));
 sky130_fd_sc_hd__nand3_1 _3985_ (.A(_2940_),
    .B(_0088_),
    .C(_0089_),
    .Y(_0106_));
 sky130_fd_sc_hd__a21o_1 _3986_ (.A1(_2940_),
    .A2(_0089_),
    .B1(_0088_),
    .X(_0107_));
 sky130_fd_sc_hd__and3_1 _3987_ (.A(_0105_),
    .B(_0106_),
    .C(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__o21ba_1 _3988_ (.A1(_2934_),
    .A2(_2937_),
    .B1_N(_2935_),
    .X(_0109_));
 sky130_fd_sc_hd__o21ba_1 _3989_ (.A1(_0090_),
    .A2(_0108_),
    .B1_N(_0109_),
    .X(_0110_));
 sky130_fd_sc_hd__or3b_1 _3990_ (.A(_0090_),
    .B(_0108_),
    .C_N(_0109_),
    .X(_0111_));
 sky130_fd_sc_hd__and2b_1 _3991_ (.A_N(_0110_),
    .B(_0111_),
    .X(_0112_));
 sky130_fd_sc_hd__a31o_2 _3992_ (.A1(_0079_),
    .A2(_2544_),
    .A3(_0112_),
    .B1(_0110_),
    .X(_0113_));
 sky130_fd_sc_hd__xor2_2 _3993_ (.A(_3086_),
    .B(_0074_),
    .X(_0114_));
 sky130_fd_sc_hd__nand2_1 _3994_ (.A(\B[2][7] ),
    .B(_2544_),
    .Y(_0115_));
 sky130_fd_sc_hd__xor2_2 _3995_ (.A(_0112_),
    .B(_0115_),
    .X(_0116_));
 sky130_fd_sc_hd__xnor2_1 _3996_ (.A(_3089_),
    .B(_0071_),
    .Y(_0117_));
 sky130_fd_sc_hd__a21oi_1 _3997_ (.A1(_0106_),
    .A2(_0107_),
    .B1(_0105_),
    .Y(_0118_));
 sky130_fd_sc_hd__nor2_1 _3998_ (.A(_0108_),
    .B(_0118_),
    .Y(_0119_));
 sky130_fd_sc_hd__or3_1 _3999_ (.A(_0069_),
    .B(_3093_),
    .C(_0068_),
    .X(_0120_));
 sky130_fd_sc_hd__o21ai_2 _4000_ (.A1(_0069_),
    .A2(_0068_),
    .B1(_3093_),
    .Y(_0121_));
 sky130_fd_sc_hd__nand3_1 _4001_ (.A(_0066_),
    .B(_3097_),
    .C(_0065_),
    .Y(_0122_));
 sky130_fd_sc_hd__a21o_1 _4002_ (.A1(_0066_),
    .A2(_0065_),
    .B1(_3097_),
    .X(_0123_));
 sky130_fd_sc_hd__xor2_1 _4003_ (.A(_0081_),
    .B(_0083_),
    .X(_0124_));
 sky130_fd_sc_hd__or3_1 _4004_ (.A(_3102_),
    .B(_3100_),
    .C(_3101_),
    .X(_0125_));
 sky130_fd_sc_hd__o21ai_1 _4005_ (.A1(_3102_),
    .A2(_3101_),
    .B1(_3100_),
    .Y(_0126_));
 sky130_fd_sc_hd__nand2_1 _4006_ (.A(_3014_),
    .B(_0960_),
    .Y(_0127_));
 sky130_fd_sc_hd__a22oi_2 _4007_ (.A1(\B[0][1] ),
    .A2(_0905_),
    .B1(_2238_),
    .B2(_3046_),
    .Y(_0128_));
 sky130_fd_sc_hd__and4_1 _4008_ (.A(\B[0][0] ),
    .B(\B[0][1] ),
    .C(\A[2][3] ),
    .D(\A[2][4] ),
    .X(_0129_));
 sky130_fd_sc_hd__o21bai_1 _4009_ (.A1(_0127_),
    .A2(_0128_),
    .B1_N(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__a21o_1 _4010_ (.A1(_0125_),
    .A2(_0126_),
    .B1(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__nand3_1 _4011_ (.A(_0125_),
    .B(_0126_),
    .C(_0130_),
    .Y(_0132_));
 sky130_fd_sc_hd__a21bo_1 _4012_ (.A1(_0124_),
    .A2(_0131_),
    .B1_N(_0132_),
    .X(_0133_));
 sky130_fd_sc_hd__and3_1 _4013_ (.A(_0122_),
    .B(_0123_),
    .C(_0133_),
    .X(_0134_));
 sky130_fd_sc_hd__nand3_1 _4014_ (.A(_0122_),
    .B(_0123_),
    .C(_0133_),
    .Y(_0135_));
 sky130_fd_sc_hd__nor3_1 _4015_ (.A(_0080_),
    .B(_0084_),
    .C(_0087_),
    .Y(_0136_));
 sky130_fd_sc_hd__nor2_1 _4016_ (.A(_0088_),
    .B(_0136_),
    .Y(_0137_));
 sky130_fd_sc_hd__a21o_1 _4017_ (.A1(_0122_),
    .A2(_0123_),
    .B1(_0133_),
    .X(_0138_));
 sky130_fd_sc_hd__and3_1 _4018_ (.A(_0135_),
    .B(_0137_),
    .C(_0138_),
    .X(_0139_));
 sky130_fd_sc_hd__a211o_2 _4019_ (.A1(_0120_),
    .A2(_0121_),
    .B1(_0134_),
    .C1(_0139_),
    .X(_0140_));
 sky130_fd_sc_hd__o211ai_4 _4020_ (.A1(_0134_),
    .A2(_0139_),
    .B1(_0120_),
    .C1(_0121_),
    .Y(_0141_));
 sky130_fd_sc_hd__a21boi_1 _4021_ (.A1(_0119_),
    .A2(_0140_),
    .B1_N(_0141_),
    .Y(_0142_));
 sky130_fd_sc_hd__xnor2_1 _4022_ (.A(_0117_),
    .B(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__nor2_1 _4023_ (.A(_0117_),
    .B(_0142_),
    .Y(_0144_));
 sky130_fd_sc_hd__o21ba_1 _4024_ (.A1(_0116_),
    .A2(_0143_),
    .B1_N(_0144_),
    .X(_0145_));
 sky130_fd_sc_hd__xnor2_2 _4025_ (.A(_0114_),
    .B(_0145_),
    .Y(_0146_));
 sky130_fd_sc_hd__and2b_1 _4026_ (.A_N(_0145_),
    .B(_0114_),
    .X(_0147_));
 sky130_fd_sc_hd__a21oi_4 _4027_ (.A1(_0113_),
    .A2(_0146_),
    .B1(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__xnor2_1 _4028_ (.A(_0078_),
    .B(_0148_),
    .Y(_0149_));
 sky130_fd_sc_hd__xnor2_2 _4029_ (.A(_0113_),
    .B(_0146_),
    .Y(_0150_));
 sky130_fd_sc_hd__xnor2_2 _4030_ (.A(_0116_),
    .B(_0143_),
    .Y(_0151_));
 sky130_fd_sc_hd__clkbuf_4 _4031_ (.A(_2895_),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_4 _4032_ (.A(_2896_),
    .X(_0153_));
 sky130_fd_sc_hd__and4_1 _4033_ (.A(_0762_),
    .B(_0883_),
    .C(_0152_),
    .D(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__and3_1 _4034_ (.A(_1740_),
    .B(_0085_),
    .C(_0154_),
    .X(_0155_));
 sky130_fd_sc_hd__a21o_1 _4035_ (.A1(_0097_),
    .A2(_0103_),
    .B1(_0102_),
    .X(_0156_));
 sky130_fd_sc_hd__and3_1 _4036_ (.A(_0104_),
    .B(_0155_),
    .C(_0156_),
    .X(_0157_));
 sky130_fd_sc_hd__and4_1 _4037_ (.A(_2916_),
    .B(\A[3][0] ),
    .C(_1598_),
    .D(_2917_),
    .X(_0158_));
 sky130_fd_sc_hd__clkbuf_4 _4038_ (.A(\B[2][5] ),
    .X(_0159_));
 sky130_fd_sc_hd__clkbuf_4 _4039_ (.A(_2917_),
    .X(_0160_));
 sky130_fd_sc_hd__a22oi_1 _4040_ (.A1(_0159_),
    .A2(_2568_),
    .B1(_1609_),
    .B2(_0160_),
    .Y(_0161_));
 sky130_fd_sc_hd__or2_1 _4041_ (.A(_0158_),
    .B(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__or3_1 _4042_ (.A(_0095_),
    .B(_0093_),
    .C(_0094_),
    .X(_0163_));
 sky130_fd_sc_hd__o21ai_1 _4043_ (.A1(_0095_),
    .A2(_0094_),
    .B1(_0093_),
    .Y(_0164_));
 sky130_fd_sc_hd__a22o_1 _4044_ (.A1(_2905_),
    .A2(_2559_),
    .B1(\A[3][3] ),
    .B2(_2903_),
    .X(_0165_));
 sky130_fd_sc_hd__and4_1 _4045_ (.A(_2903_),
    .B(\B[2][2] ),
    .C(_2559_),
    .D(\A[3][3] ),
    .X(_0166_));
 sky130_fd_sc_hd__a31o_1 _4046_ (.A1(_1598_),
    .A2(\B[2][3] ),
    .A3(_0165_),
    .B1(_0166_),
    .X(_0167_));
 sky130_fd_sc_hd__a21oi_1 _4047_ (.A1(_0163_),
    .A2(_0164_),
    .B1(_0167_),
    .Y(_0168_));
 sky130_fd_sc_hd__and3_1 _4048_ (.A(_0163_),
    .B(_0164_),
    .C(_0167_),
    .X(_0169_));
 sky130_fd_sc_hd__o21ba_1 _4049_ (.A1(_0162_),
    .A2(_0168_),
    .B1_N(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__inv_2 _4050_ (.A(_0170_),
    .Y(_0171_));
 sky130_fd_sc_hd__nand3_1 _4051_ (.A(_0104_),
    .B(_0155_),
    .C(_0156_),
    .Y(_0172_));
 sky130_fd_sc_hd__a21o_1 _4052_ (.A1(_0104_),
    .A2(_0156_),
    .B1(_0155_),
    .X(_0173_));
 sky130_fd_sc_hd__and3_1 _4053_ (.A(_0171_),
    .B(_0172_),
    .C(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__o21ba_1 _4054_ (.A1(_0098_),
    .A2(_0101_),
    .B1_N(_0099_),
    .X(_0175_));
 sky130_fd_sc_hd__o21ba_1 _4055_ (.A1(_0157_),
    .A2(_0174_),
    .B1_N(_0175_),
    .X(_0176_));
 sky130_fd_sc_hd__or3b_1 _4056_ (.A(_0157_),
    .B(_0174_),
    .C_N(_0175_),
    .X(_0177_));
 sky130_fd_sc_hd__and2b_1 _4057_ (.A_N(_0176_),
    .B(_0177_),
    .X(_0178_));
 sky130_fd_sc_hd__nand2_1 _4058_ (.A(_2886_),
    .B(_2717_),
    .Y(_0179_));
 sky130_fd_sc_hd__xnor2_1 _4059_ (.A(_0178_),
    .B(_0179_),
    .Y(_0180_));
 sky130_fd_sc_hd__and3_1 _4060_ (.A(_0141_),
    .B(_0119_),
    .C(_0140_),
    .X(_0181_));
 sky130_fd_sc_hd__a21oi_2 _4061_ (.A1(_0141_),
    .A2(_0140_),
    .B1(_0119_),
    .Y(_0182_));
 sky130_fd_sc_hd__nand3_1 _4062_ (.A(_0132_),
    .B(_0124_),
    .C(_0131_),
    .Y(_0183_));
 sky130_fd_sc_hd__a21o_1 _4063_ (.A1(_0132_),
    .A2(_0131_),
    .B1(_0124_),
    .X(_0184_));
 sky130_fd_sc_hd__buf_4 _4064_ (.A(_2895_),
    .X(_0185_));
 sky130_fd_sc_hd__buf_4 _4065_ (.A(_0153_),
    .X(_0186_));
 sky130_fd_sc_hd__a22oi_1 _4066_ (.A1(_0883_),
    .A2(_0185_),
    .B1(_0186_),
    .B2(_0773_),
    .Y(_0187_));
 sky130_fd_sc_hd__nor2_1 _4067_ (.A(_0154_),
    .B(_0187_),
    .Y(_0188_));
 sky130_fd_sc_hd__or3_1 _4068_ (.A(_0129_),
    .B(_0127_),
    .C(_0128_),
    .X(_0189_));
 sky130_fd_sc_hd__o21ai_1 _4069_ (.A1(_0129_),
    .A2(_0128_),
    .B1(_0127_),
    .Y(_0190_));
 sky130_fd_sc_hd__nand2_1 _4070_ (.A(_0817_),
    .B(_3014_),
    .Y(_0191_));
 sky130_fd_sc_hd__a22oi_2 _4071_ (.A1(_3015_),
    .A2(_0960_),
    .B1(_1004_),
    .B2(_3046_),
    .Y(_0192_));
 sky130_fd_sc_hd__and4_1 _4072_ (.A(_3046_),
    .B(\B[0][1] ),
    .C(_0960_),
    .D(_0905_),
    .X(_0193_));
 sky130_fd_sc_hd__o21bai_1 _4073_ (.A1(_0191_),
    .A2(_0192_),
    .B1_N(_0193_),
    .Y(_0194_));
 sky130_fd_sc_hd__a21o_1 _4074_ (.A1(_0189_),
    .A2(_0190_),
    .B1(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__nand3_1 _4075_ (.A(_0189_),
    .B(_0190_),
    .C(_0194_),
    .Y(_0196_));
 sky130_fd_sc_hd__a21bo_1 _4076_ (.A1(_0188_),
    .A2(_0195_),
    .B1_N(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__and3_2 _4077_ (.A(_0183_),
    .B(_0184_),
    .C(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__a21oi_1 _4078_ (.A1(_2676_),
    .A2(_0085_),
    .B1(_0154_),
    .Y(_0199_));
 sky130_fd_sc_hd__or2_1 _4079_ (.A(_0155_),
    .B(_0199_),
    .X(_0200_));
 sky130_fd_sc_hd__a21oi_2 _4080_ (.A1(_0183_),
    .A2(_0184_),
    .B1(_0197_),
    .Y(_0201_));
 sky130_fd_sc_hd__nor3_4 _4081_ (.A(_0198_),
    .B(_0200_),
    .C(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__nand3_2 _4082_ (.A(_0135_),
    .B(_0137_),
    .C(_0138_),
    .Y(_0203_));
 sky130_fd_sc_hd__a21o_1 _4083_ (.A1(_0135_),
    .A2(_0138_),
    .B1(_0137_),
    .X(_0204_));
 sky130_fd_sc_hd__o211a_2 _4084_ (.A1(_0198_),
    .A2(_0202_),
    .B1(_0203_),
    .C1(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__inv_2 _4085_ (.A(_0205_),
    .Y(_0206_));
 sky130_fd_sc_hd__a21oi_1 _4086_ (.A1(_0172_),
    .A2(_0173_),
    .B1(_0171_),
    .Y(_0207_));
 sky130_fd_sc_hd__or2_1 _4087_ (.A(_0174_),
    .B(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__a211oi_4 _4088_ (.A1(_0203_),
    .A2(_0204_),
    .B1(_0198_),
    .C1(_0202_),
    .Y(_0209_));
 sky130_fd_sc_hd__or3_1 _4089_ (.A(_0205_),
    .B(_0208_),
    .C(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__o211ai_2 _4090_ (.A1(_0181_),
    .A2(_0182_),
    .B1(_0206_),
    .C1(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__a211o_1 _4091_ (.A1(_0206_),
    .A2(_0210_),
    .B1(_0181_),
    .C1(_0182_),
    .X(_0212_));
 sky130_fd_sc_hd__a21bo_1 _4092_ (.A1(_0180_),
    .A2(_0211_),
    .B1_N(_0212_),
    .X(_0213_));
 sky130_fd_sc_hd__or2b_1 _4093_ (.A(_0151_),
    .B_N(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__a31o_1 _4094_ (.A1(_2886_),
    .A2(_2717_),
    .A3(_0178_),
    .B1(_0176_),
    .X(_0215_));
 sky130_fd_sc_hd__xnor2_1 _4095_ (.A(_0151_),
    .B(_0213_),
    .Y(_0216_));
 sky130_fd_sc_hd__nand2_1 _4096_ (.A(_0215_),
    .B(_0216_),
    .Y(_0217_));
 sky130_fd_sc_hd__and3_1 _4097_ (.A(_0150_),
    .B(_0214_),
    .C(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__and4_1 _4098_ (.A(_2903_),
    .B(\A[3][1] ),
    .C(_2905_),
    .D(_2559_),
    .X(_0219_));
 sky130_fd_sc_hd__clkbuf_4 _4099_ (.A(\B[2][2] ),
    .X(_0220_));
 sky130_fd_sc_hd__clkbuf_4 _4100_ (.A(\B[2][1] ),
    .X(_0221_));
 sky130_fd_sc_hd__a22oi_1 _4101_ (.A1(_1598_),
    .A2(_0220_),
    .B1(_0707_),
    .B2(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__and4bb_1 _4102_ (.A_N(_0219_),
    .B_N(_0222_),
    .C(_2568_),
    .D(_3001_),
    .X(_0223_));
 sky130_fd_sc_hd__nor2_1 _4103_ (.A(_0219_),
    .B(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__nand2_1 _4104_ (.A(_1609_),
    .B(_3001_),
    .Y(_0225_));
 sky130_fd_sc_hd__and2b_1 _4105_ (.A_N(_0166_),
    .B(_0165_),
    .X(_0226_));
 sky130_fd_sc_hd__xnor2_1 _4106_ (.A(_0225_),
    .B(_0226_),
    .Y(_0227_));
 sky130_fd_sc_hd__and2b_1 _4107_ (.A_N(_0224_),
    .B(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__buf_4 _4108_ (.A(_2917_),
    .X(_0229_));
 sky130_fd_sc_hd__xnor2_1 _4109_ (.A(_0227_),
    .B(_0224_),
    .Y(_0230_));
 sky130_fd_sc_hd__and3_1 _4110_ (.A(_2629_),
    .B(_0229_),
    .C(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__nor2_1 _4111_ (.A(_0169_),
    .B(_0168_),
    .Y(_0232_));
 sky130_fd_sc_hd__xnor2_1 _4112_ (.A(_0162_),
    .B(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__o21a_1 _4113_ (.A1(_0228_),
    .A2(_0231_),
    .B1(_0233_),
    .X(_0234_));
 sky130_fd_sc_hd__and2_1 _4114_ (.A(_0158_),
    .B(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__nand3_1 _4115_ (.A(_0196_),
    .B(_0188_),
    .C(_0195_),
    .Y(_0236_));
 sky130_fd_sc_hd__a21o_1 _4116_ (.A1(_0196_),
    .A2(_0195_),
    .B1(_0188_),
    .X(_0237_));
 sky130_fd_sc_hd__nand2_1 _4117_ (.A(_2550_),
    .B(_0185_),
    .Y(_0238_));
 sky130_fd_sc_hd__or3_1 _4118_ (.A(_0193_),
    .B(_0191_),
    .C(_0192_),
    .X(_0239_));
 sky130_fd_sc_hd__o21ai_1 _4119_ (.A1(_0193_),
    .A2(_0192_),
    .B1(_0191_),
    .Y(_0240_));
 sky130_fd_sc_hd__buf_4 _4120_ (.A(_3014_),
    .X(_0241_));
 sky130_fd_sc_hd__a22o_1 _4121_ (.A1(_3015_),
    .A2(_0872_),
    .B1(_0993_),
    .B2(_3046_),
    .X(_0242_));
 sky130_fd_sc_hd__and4_1 _4122_ (.A(_3046_),
    .B(_3015_),
    .C(_0872_),
    .D(_0993_),
    .X(_0243_));
 sky130_fd_sc_hd__a31o_1 _4123_ (.A1(_0762_),
    .A2(_0241_),
    .A3(_0242_),
    .B1(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__a21oi_2 _4124_ (.A1(_0239_),
    .A2(_0240_),
    .B1(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__and3_1 _4125_ (.A(_0239_),
    .B(_0240_),
    .C(_0244_),
    .X(_0246_));
 sky130_fd_sc_hd__o21bai_2 _4126_ (.A1(_0238_),
    .A2(_0245_),
    .B1_N(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__nand3_4 _4127_ (.A(_0236_),
    .B(_0237_),
    .C(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__buf_4 _4128_ (.A(_0085_),
    .X(_0249_));
 sky130_fd_sc_hd__a21o_1 _4129_ (.A1(_0236_),
    .A2(_0237_),
    .B1(_0247_),
    .X(_0250_));
 sky130_fd_sc_hd__nand4_4 _4130_ (.A(_0249_),
    .B(_2668_),
    .C(_0248_),
    .D(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__o21a_1 _4131_ (.A1(_0198_),
    .A2(_0201_),
    .B1(_0200_),
    .X(_0252_));
 sky130_fd_sc_hd__a211oi_4 _4132_ (.A1(_0248_),
    .A2(_0251_),
    .B1(_0202_),
    .C1(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__inv_2 _4133_ (.A(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__o211a_1 _4134_ (.A1(_0202_),
    .A2(_0252_),
    .B1(_0248_),
    .C1(_0251_),
    .X(_0255_));
 sky130_fd_sc_hd__nor3_1 _4135_ (.A(_0228_),
    .B(_0231_),
    .C(_0233_),
    .Y(_0256_));
 sky130_fd_sc_hd__nor2_1 _4136_ (.A(_0234_),
    .B(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__or3b_4 _4137_ (.A(_0253_),
    .B(_0255_),
    .C_N(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__nor3_2 _4138_ (.A(_0205_),
    .B(_0208_),
    .C(_0209_),
    .Y(_0259_));
 sky130_fd_sc_hd__o21a_1 _4139_ (.A1(_0205_),
    .A2(_0209_),
    .B1(_0208_),
    .X(_0260_));
 sky130_fd_sc_hd__a211oi_4 _4140_ (.A1(_0254_),
    .A2(_0258_),
    .B1(_0259_),
    .C1(_0260_),
    .Y(_0261_));
 sky130_fd_sc_hd__nor2_1 _4141_ (.A(_0158_),
    .B(_0234_),
    .Y(_0262_));
 sky130_fd_sc_hd__or2_1 _4142_ (.A(_0235_),
    .B(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__o211a_1 _4143_ (.A1(_0259_),
    .A2(_0260_),
    .B1(_0254_),
    .C1(_0258_),
    .X(_0264_));
 sky130_fd_sc_hd__nor3_2 _4144_ (.A(_0261_),
    .B(_0263_),
    .C(_0264_),
    .Y(_0265_));
 sky130_fd_sc_hd__nand3_1 _4145_ (.A(_0212_),
    .B(_0180_),
    .C(_0211_),
    .Y(_0266_));
 sky130_fd_sc_hd__a21o_1 _4146_ (.A1(_0212_),
    .A2(_0211_),
    .B1(_0180_),
    .X(_0267_));
 sky130_fd_sc_hd__o211ai_2 _4147_ (.A1(_0261_),
    .A2(_0265_),
    .B1(_0266_),
    .C1(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__a211o_1 _4148_ (.A1(_0266_),
    .A2(_0267_),
    .B1(_0261_),
    .C1(_0265_),
    .X(_0269_));
 sky130_fd_sc_hd__nand3_1 _4149_ (.A(_0235_),
    .B(_0268_),
    .C(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__a21o_1 _4150_ (.A1(_0268_),
    .A2(_0269_),
    .B1(_0235_),
    .X(_0271_));
 sky130_fd_sc_hd__a22o_1 _4151_ (.A1(_0249_),
    .A2(_2668_),
    .B1(_0248_),
    .B2(_0250_),
    .X(_0272_));
 sky130_fd_sc_hd__and2_1 _4152_ (.A(_0249_),
    .B(_1532_),
    .X(_0273_));
 sky130_fd_sc_hd__or3_1 _4153_ (.A(_0238_),
    .B(_0246_),
    .C(_0245_),
    .X(_0274_));
 sky130_fd_sc_hd__o21ai_2 _4154_ (.A1(_0246_),
    .A2(_0245_),
    .B1(_0238_),
    .Y(_0275_));
 sky130_fd_sc_hd__nand2_1 _4155_ (.A(_0773_),
    .B(_0241_),
    .Y(_0276_));
 sky130_fd_sc_hd__and2b_1 _4156_ (.A_N(_0243_),
    .B(_0242_),
    .X(_0277_));
 sky130_fd_sc_hd__xnor2_2 _4157_ (.A(_0276_),
    .B(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__clkbuf_4 _4158_ (.A(\B[0][0] ),
    .X(_0279_));
 sky130_fd_sc_hd__buf_4 _4159_ (.A(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__buf_2 _4160_ (.A(\B[0][1] ),
    .X(_0281_));
 sky130_fd_sc_hd__buf_4 _4161_ (.A(_0281_),
    .X(_0282_));
 sky130_fd_sc_hd__and4_1 _4162_ (.A(_0280_),
    .B(_0773_),
    .C(_0282_),
    .D(_0883_),
    .X(_0283_));
 sky130_fd_sc_hd__and2_1 _4163_ (.A(_0278_),
    .B(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__a21o_1 _4164_ (.A1(_0274_),
    .A2(_0275_),
    .B1(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__nand3_1 _4165_ (.A(_0274_),
    .B(_0275_),
    .C(_0284_),
    .Y(_0286_));
 sky130_fd_sc_hd__a21bo_1 _4166_ (.A1(_0273_),
    .A2(_0285_),
    .B1_N(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__and3_2 _4167_ (.A(_0251_),
    .B(_0272_),
    .C(_0287_),
    .X(_0288_));
 sky130_fd_sc_hd__nand2_1 _4168_ (.A(_2629_),
    .B(_0229_),
    .Y(_0289_));
 sky130_fd_sc_hd__xnor2_1 _4169_ (.A(_0289_),
    .B(_0230_),
    .Y(_0290_));
 sky130_fd_sc_hd__o2bb2a_1 _4170_ (.A1_N(_2568_),
    .A2_N(_3002_),
    .B1(_0219_),
    .B2(_0222_),
    .X(_0291_));
 sky130_fd_sc_hd__nor2_1 _4171_ (.A(_0223_),
    .B(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__clkbuf_4 _4172_ (.A(_2903_),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_4 _4173_ (.A(_2905_),
    .X(_0294_));
 sky130_fd_sc_hd__and4_1 _4174_ (.A(_2629_),
    .B(_0293_),
    .C(_1609_),
    .D(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__and2_1 _4175_ (.A(_0292_),
    .B(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__and2_1 _4176_ (.A(_0290_),
    .B(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__nor2_1 _4177_ (.A(_0290_),
    .B(_0296_),
    .Y(_0298_));
 sky130_fd_sc_hd__or2_1 _4178_ (.A(_0297_),
    .B(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__a21oi_2 _4179_ (.A1(_0251_),
    .A2(_0272_),
    .B1(_0287_),
    .Y(_0300_));
 sky130_fd_sc_hd__nor3_1 _4180_ (.A(_0288_),
    .B(_0299_),
    .C(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__o21bai_1 _4181_ (.A1(_0253_),
    .A2(_0255_),
    .B1_N(_0257_),
    .Y(_0302_));
 sky130_fd_sc_hd__o211ai_2 _4182_ (.A1(_0288_),
    .A2(_0301_),
    .B1(_0258_),
    .C1(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__a211o_1 _4183_ (.A1(_0258_),
    .A2(_0302_),
    .B1(_0288_),
    .C1(_0301_),
    .X(_0304_));
 sky130_fd_sc_hd__nand3_1 _4184_ (.A(_0297_),
    .B(_0303_),
    .C(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__o21a_1 _4185_ (.A1(_0261_),
    .A2(_0264_),
    .B1(_0263_),
    .X(_0306_));
 sky130_fd_sc_hd__a211oi_2 _4186_ (.A1(_0303_),
    .A2(_0305_),
    .B1(_0306_),
    .C1(_0265_),
    .Y(_0307_));
 sky130_fd_sc_hd__a21oi_1 _4187_ (.A1(_0270_),
    .A2(_0271_),
    .B1(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__or3_1 _4188_ (.A(_0288_),
    .B(_0299_),
    .C(_0300_),
    .X(_0309_));
 sky130_fd_sc_hd__o21ai_1 _4189_ (.A1(_0288_),
    .A2(_0300_),
    .B1(_0299_),
    .Y(_0310_));
 sky130_fd_sc_hd__nand3_1 _4190_ (.A(_0286_),
    .B(_0273_),
    .C(_0285_),
    .Y(_0311_));
 sky130_fd_sc_hd__a21o_1 _4191_ (.A1(_0286_),
    .A2(_0285_),
    .B1(_0273_),
    .X(_0312_));
 sky130_fd_sc_hd__inv_2 _4192_ (.A(_0283_),
    .Y(_0313_));
 sky130_fd_sc_hd__xnor2_1 _4193_ (.A(_0278_),
    .B(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__and3_1 _4194_ (.A(_0249_),
    .B(_0718_),
    .C(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__a21o_1 _4195_ (.A1(_0311_),
    .A2(_0312_),
    .B1(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__nor2_1 _4196_ (.A(_0292_),
    .B(_0295_),
    .Y(_0317_));
 sky130_fd_sc_hd__nor2_1 _4197_ (.A(_0296_),
    .B(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__nand3_1 _4198_ (.A(_0311_),
    .B(_0312_),
    .C(_0315_),
    .Y(_0319_));
 sky130_fd_sc_hd__a21bo_1 _4199_ (.A1(_0316_),
    .A2(_0318_),
    .B1_N(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__and3_1 _4200_ (.A(_0309_),
    .B(_0310_),
    .C(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__a21o_1 _4201_ (.A1(_0309_),
    .A2(_0310_),
    .B1(_0320_),
    .X(_0322_));
 sky130_fd_sc_hd__nand3_1 _4202_ (.A(_0319_),
    .B(_0316_),
    .C(_0318_),
    .Y(_0323_));
 sky130_fd_sc_hd__a21o_1 _4203_ (.A1(_0319_),
    .A2(_0316_),
    .B1(_0318_),
    .X(_0324_));
 sky130_fd_sc_hd__nand2_1 _4204_ (.A(_0249_),
    .B(_0718_),
    .Y(_0325_));
 sky130_fd_sc_hd__xnor2_1 _4205_ (.A(_0314_),
    .B(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__a22o_1 _4206_ (.A1(_2550_),
    .A2(_0282_),
    .B1(_0883_),
    .B2(_0280_),
    .X(_0327_));
 sky130_fd_sc_hd__and4_1 _4207_ (.A(_0249_),
    .B(_1609_),
    .C(_0313_),
    .D(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__xnor2_1 _4208_ (.A(_0326_),
    .B(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__a22oi_1 _4209_ (.A1(_0293_),
    .A2(_2544_),
    .B1(_0294_),
    .B2(_2629_),
    .Y(_0330_));
 sky130_fd_sc_hd__or2_1 _4210_ (.A(_0295_),
    .B(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__nor2_1 _4211_ (.A(_0329_),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__a21o_1 _4212_ (.A1(_0326_),
    .A2(_0328_),
    .B1(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__and3_1 _4213_ (.A(_0323_),
    .B(_0324_),
    .C(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__and3b_1 _4214_ (.A_N(_0321_),
    .B(_0322_),
    .C(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__a21o_1 _4215_ (.A1(_0303_),
    .A2(_0304_),
    .B1(_0297_),
    .X(_0336_));
 sky130_fd_sc_hd__and2_1 _4216_ (.A(_0305_),
    .B(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__and2b_1 _4217_ (.A_N(_0321_),
    .B(_0322_),
    .X(_0338_));
 sky130_fd_sc_hd__a21oi_1 _4218_ (.A1(_0323_),
    .A2(_0324_),
    .B1(_0333_),
    .Y(_0339_));
 sky130_fd_sc_hd__and2_1 _4219_ (.A(_0329_),
    .B(_0331_),
    .X(_0340_));
 sky130_fd_sc_hd__nor2_1 _4220_ (.A(_0332_),
    .B(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__clkbuf_4 _4221_ (.A(_0249_),
    .X(_0342_));
 sky130_fd_sc_hd__a22oi_1 _4222_ (.A1(_0342_),
    .A2(_2544_),
    .B1(_0313_),
    .B2(_0327_),
    .Y(_0343_));
 sky130_fd_sc_hd__nor2_1 _4223_ (.A(_0328_),
    .B(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__and4_1 _4224_ (.A(_0280_),
    .B(_0342_),
    .C(_2550_),
    .D(_2717_),
    .X(_0345_));
 sky130_fd_sc_hd__nand2_1 _4225_ (.A(_2717_),
    .B(_0293_),
    .Y(_0346_));
 sky130_fd_sc_hd__xnor2_1 _4226_ (.A(_0344_),
    .B(_0345_),
    .Y(_0347_));
 sky130_fd_sc_hd__nor2_1 _4227_ (.A(_0346_),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__a21o_1 _4228_ (.A1(_0344_),
    .A2(_0345_),
    .B1(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__nand2_1 _4229_ (.A(_0341_),
    .B(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__nor3_1 _4230_ (.A(_0334_),
    .B(_0339_),
    .C(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__and2_1 _4231_ (.A(_0338_),
    .B(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__nor2_1 _4232_ (.A(_0321_),
    .B(_0335_),
    .Y(_0353_));
 sky130_fd_sc_hd__xnor2_1 _4233_ (.A(_0337_),
    .B(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__a22oi_2 _4234_ (.A1(_0335_),
    .A2(_0337_),
    .B1(_0352_),
    .B2(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__o211a_1 _4235_ (.A1(_0265_),
    .A2(_0306_),
    .B1(_0305_),
    .C1(_0303_),
    .X(_0356_));
 sky130_fd_sc_hd__and4bb_1 _4236_ (.A_N(_0307_),
    .B_N(_0356_),
    .C(_0337_),
    .D(_0321_),
    .X(_0357_));
 sky130_fd_sc_hd__o2bb2a_1 _4237_ (.A1_N(_0321_),
    .A2_N(_0337_),
    .B1(_0356_),
    .B2(_0307_),
    .X(_0358_));
 sky130_fd_sc_hd__or2_1 _4238_ (.A(_0357_),
    .B(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__o211ai_1 _4239_ (.A1(_0307_),
    .A2(_0357_),
    .B1(_0270_),
    .C1(_0271_),
    .Y(_0360_));
 sky130_fd_sc_hd__o31a_1 _4240_ (.A1(_0308_),
    .A2(_0355_),
    .A3(_0359_),
    .B1(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__or2_1 _4241_ (.A(_0215_),
    .B(_0216_),
    .X(_0362_));
 sky130_fd_sc_hd__and2_1 _4242_ (.A(_0217_),
    .B(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__and2_1 _4243_ (.A(_0268_),
    .B(_0270_),
    .X(_0364_));
 sky130_fd_sc_hd__xor2_2 _4244_ (.A(_0363_),
    .B(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__or2b_1 _4245_ (.A(_0364_),
    .B_N(_0363_),
    .X(_0366_));
 sky130_fd_sc_hd__o21ai_1 _4246_ (.A1(_0361_),
    .A2(_0365_),
    .B1(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__a21o_1 _4247_ (.A1(_0214_),
    .A2(_0217_),
    .B1(_0150_),
    .X(_0368_));
 sky130_fd_sc_hd__and2b_1 _4248_ (.A_N(_0367_),
    .B(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__or3_1 _4249_ (.A(_0149_),
    .B(_0218_),
    .C(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__o21ai_1 _4250_ (.A1(_0078_),
    .A2(_0148_),
    .B1(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__nor2_1 _4251_ (.A(_3084_),
    .B(_0076_),
    .Y(_0372_));
 sky130_fd_sc_hd__a21oi_2 _4252_ (.A1(_2947_),
    .A2(_0077_),
    .B1(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__a31o_2 _4253_ (.A1(_0079_),
    .A2(_1532_),
    .A3(_2978_),
    .B1(_2976_),
    .X(_0374_));
 sky130_fd_sc_hd__nor2_1 _4254_ (.A(_3059_),
    .B(_3082_),
    .Y(_0375_));
 sky130_fd_sc_hd__a21o_1 _4255_ (.A1(_2980_),
    .A2(_3083_),
    .B1(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__nand2_1 _4256_ (.A(_2886_),
    .B(_2668_),
    .Y(_0377_));
 sky130_fd_sc_hd__buf_4 _4257_ (.A(_0159_),
    .X(_0378_));
 sky130_fd_sc_hd__and4_1 _4258_ (.A(_0378_),
    .B(_2551_),
    .C(_2676_),
    .D(_0229_),
    .X(_0379_));
 sky130_fd_sc_hd__or2_1 _4259_ (.A(_0379_),
    .B(_2999_),
    .X(_0380_));
 sky130_fd_sc_hd__a21oi_4 _4260_ (.A1(_2984_),
    .A2(_3006_),
    .B1(_3005_),
    .Y(_0381_));
 sky130_fd_sc_hd__xnor2_2 _4261_ (.A(_0380_),
    .B(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__xnor2_2 _4262_ (.A(_0377_),
    .B(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__and2_1 _4263_ (.A(_3038_),
    .B(_3057_),
    .X(_0384_));
 sky130_fd_sc_hd__a21oi_2 _4264_ (.A1(_3008_),
    .A2(_3058_),
    .B1(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__a21oi_2 _4265_ (.A1(_3000_),
    .A2(_3003_),
    .B1(_2982_),
    .Y(_0386_));
 sky130_fd_sc_hd__and2b_1 _4266_ (.A_N(_3033_),
    .B(_3029_),
    .X(_0387_));
 sky130_fd_sc_hd__buf_4 _4267_ (.A(_2921_),
    .X(_0388_));
 sky130_fd_sc_hd__nand2_1 _4268_ (.A(_0388_),
    .B(_2676_),
    .Y(_0389_));
 sky130_fd_sc_hd__a22oi_1 _4269_ (.A1(_0378_),
    .A2(_2551_),
    .B1(_0229_),
    .B2(_0806_),
    .Y(_0390_));
 sky130_fd_sc_hd__and4_1 _4270_ (.A(_0378_),
    .B(_0806_),
    .C(_0751_),
    .D(_0160_),
    .X(_0391_));
 sky130_fd_sc_hd__nor2_1 _4271_ (.A(_0390_),
    .B(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__xnor2_1 _4272_ (.A(_0389_),
    .B(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__o21a_1 _4273_ (.A1(_0387_),
    .A2(_3036_),
    .B1(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__nor3_1 _4274_ (.A(_0387_),
    .B(_3036_),
    .C(_0393_),
    .Y(_0395_));
 sky130_fd_sc_hd__nor2_1 _4275_ (.A(_0394_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__xnor2_2 _4276_ (.A(_0386_),
    .B(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__a21oi_2 _4277_ (.A1(_3027_),
    .A2(_3037_),
    .B1(_3026_),
    .Y(_0398_));
 sky130_fd_sc_hd__nand2_2 _4278_ (.A(_2988_),
    .B(_2431_),
    .Y(_0399_));
 sky130_fd_sc_hd__buf_4 _4279_ (.A(_2988_),
    .X(_0400_));
 sky130_fd_sc_hd__a22o_1 _4280_ (.A1(_0400_),
    .A2(_2858_),
    .B1(_0186_),
    .B2(_2859_),
    .X(_0401_));
 sky130_fd_sc_hd__o21ai_2 _4281_ (.A1(_3021_),
    .A2(_0399_),
    .B1(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__a22o_1 _4282_ (.A1(_2888_),
    .A2(_2445_),
    .B1(_1915_),
    .B2(_2964_),
    .X(_0403_));
 sky130_fd_sc_hd__nand2_1 _4283_ (.A(_2964_),
    .B(_2218_),
    .Y(_0404_));
 sky130_fd_sc_hd__or2_1 _4284_ (.A(_3031_),
    .B(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__nand2_1 _4285_ (.A(_0403_),
    .B(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__a31o_1 _4286_ (.A1(_0400_),
    .A2(_2445_),
    .A3(_3023_),
    .B1(_3022_),
    .X(_0407_));
 sky130_fd_sc_hd__xor2_1 _4287_ (.A(_0406_),
    .B(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__xnor2_1 _4288_ (.A(_3032_),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__xnor2_2 _4289_ (.A(_0402_),
    .B(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__xnor2_2 _4290_ (.A(_0398_),
    .B(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__xnor2_2 _4291_ (.A(_0397_),
    .B(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__xor2_2 _4292_ (.A(_0385_),
    .B(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__xnor2_2 _4293_ (.A(_0383_),
    .B(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__xnor2_2 _4294_ (.A(_0376_),
    .B(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__xnor2_4 _4295_ (.A(_0374_),
    .B(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__xnor2_1 _4296_ (.A(_0373_),
    .B(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__xnor2_1 _4297_ (.A(_0371_),
    .B(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__buf_2 _4298_ (.A(\A[1][2] ),
    .X(_0419_));
 sky130_fd_sc_hd__buf_2 _4299_ (.A(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_4 _4300_ (.A(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__buf_2 _4301_ (.A(\A[1][6] ),
    .X(_0422_));
 sky130_fd_sc_hd__nand4_1 _4302_ (.A(\A[1][7] ),
    .B(_0422_),
    .C(_1136_),
    .D(_1103_),
    .Y(_0423_));
 sky130_fd_sc_hd__a22o_1 _4303_ (.A1(\A[1][7] ),
    .A2(_1092_),
    .B1(_1257_),
    .B2(_0422_),
    .X(_0424_));
 sky130_fd_sc_hd__buf_2 _4304_ (.A(\A[1][5] ),
    .X(_0425_));
 sky130_fd_sc_hd__and2_1 _4305_ (.A(_0425_),
    .B(\B[3][3] ),
    .X(_0426_));
 sky130_fd_sc_hd__nand3_1 _4306_ (.A(_0423_),
    .B(_0424_),
    .C(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__a21o_1 _4307_ (.A1(_0423_),
    .A2(_0424_),
    .B1(_0426_),
    .X(_0428_));
 sky130_fd_sc_hd__a22oi_2 _4308_ (.A1(_0422_),
    .A2(_1136_),
    .B1(_1103_),
    .B2(_0425_),
    .Y(_0429_));
 sky130_fd_sc_hd__buf_2 _4309_ (.A(\A[1][4] ),
    .X(_0430_));
 sky130_fd_sc_hd__nand2_1 _4310_ (.A(_1202_),
    .B(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__and4_1 _4311_ (.A(\A[1][6] ),
    .B(\A[1][5] ),
    .C(_1092_),
    .D(\B[3][2] ),
    .X(_0432_));
 sky130_fd_sc_hd__o21bai_1 _4312_ (.A1(_0429_),
    .A2(_0431_),
    .B1_N(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__and3_1 _4313_ (.A(_0427_),
    .B(_0428_),
    .C(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__a21oi_1 _4314_ (.A1(_0427_),
    .A2(_0428_),
    .B1(_0433_),
    .Y(_0435_));
 sky130_fd_sc_hd__buf_2 _4315_ (.A(\A[1][3] ),
    .X(_0436_));
 sky130_fd_sc_hd__a22oi_1 _4316_ (.A1(_1312_),
    .A2(_0436_),
    .B1(_0430_),
    .B2(_1334_),
    .Y(_0437_));
 sky130_fd_sc_hd__and4_1 _4317_ (.A(\B[3][5] ),
    .B(_0436_),
    .C(_0430_),
    .D(\B[3][4] ),
    .X(_0438_));
 sky130_fd_sc_hd__nor2_1 _4318_ (.A(_0437_),
    .B(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__nand2_1 _4319_ (.A(\B[3][6] ),
    .B(_0420_),
    .Y(_0440_));
 sky130_fd_sc_hd__xnor2_1 _4320_ (.A(_0439_),
    .B(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__or3b_1 _4321_ (.A(_0434_),
    .B(_0435_),
    .C_N(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_4 _4322_ (.A(_0422_),
    .X(_0443_));
 sky130_fd_sc_hd__buf_2 _4323_ (.A(\A[0][0] ),
    .X(_0444_));
 sky130_fd_sc_hd__and4_1 _4324_ (.A(_0443_),
    .B(_0729_),
    .C(_0444_),
    .D(_0784_),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_4 _4325_ (.A(\A[1][7] ),
    .X(_0446_));
 sky130_fd_sc_hd__buf_2 _4326_ (.A(\A[0][1] ),
    .X(_0447_));
 sky130_fd_sc_hd__nand4_1 _4327_ (.A(\B[1][6] ),
    .B(\B[1][7] ),
    .C(\A[0][0] ),
    .D(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__a22o_1 _4328_ (.A1(\B[1][7] ),
    .A2(\A[0][0] ),
    .B1(_0447_),
    .B2(\B[1][6] ),
    .X(_0449_));
 sky130_fd_sc_hd__nand4_1 _4329_ (.A(_0446_),
    .B(\B[3][0] ),
    .C(_0448_),
    .D(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__a22o_1 _4330_ (.A1(\A[1][7] ),
    .A2(\B[3][0] ),
    .B1(_0448_),
    .B2(_0449_),
    .X(_0451_));
 sky130_fd_sc_hd__nand2_1 _4331_ (.A(\B[1][5] ),
    .B(_0447_),
    .Y(_0452_));
 sky130_fd_sc_hd__clkbuf_4 _4332_ (.A(\A[0][3] ),
    .X(_0453_));
 sky130_fd_sc_hd__buf_2 _4333_ (.A(net53),
    .X(_0454_));
 sky130_fd_sc_hd__buf_2 _4334_ (.A(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__a22oi_1 _4335_ (.A1(_0453_),
    .A2(_0927_),
    .B1(_1026_),
    .B2(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__buf_2 _4336_ (.A(net52),
    .X(_0457_));
 sky130_fd_sc_hd__and4_1 _4337_ (.A(_0454_),
    .B(_0457_),
    .C(_1015_),
    .D(_0938_),
    .X(_0458_));
 sky130_fd_sc_hd__o21bai_1 _4338_ (.A1(_0452_),
    .A2(_0456_),
    .B1_N(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__a21o_1 _4339_ (.A1(_0450_),
    .A2(_0451_),
    .B1(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__nand3_1 _4340_ (.A(_0450_),
    .B(_0459_),
    .C(_0451_),
    .Y(_0461_));
 sky130_fd_sc_hd__a21bo_1 _4341_ (.A1(_0445_),
    .A2(_0460_),
    .B1_N(_0461_),
    .X(_0462_));
 sky130_fd_sc_hd__o21bai_1 _4342_ (.A1(_0434_),
    .A2(_0435_),
    .B1_N(_0441_),
    .Y(_0463_));
 sky130_fd_sc_hd__and3_1 _4343_ (.A(_0442_),
    .B(_0462_),
    .C(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__or3_1 _4344_ (.A(_0432_),
    .B(_0429_),
    .C(_0431_),
    .X(_0465_));
 sky130_fd_sc_hd__o21ai_1 _4345_ (.A1(_0432_),
    .A2(_0429_),
    .B1(_0431_),
    .Y(_0466_));
 sky130_fd_sc_hd__a22oi_2 _4346_ (.A1(_0425_),
    .A2(_1136_),
    .B1(_1103_),
    .B2(_0430_),
    .Y(_0467_));
 sky130_fd_sc_hd__nand2_1 _4347_ (.A(_0436_),
    .B(_1202_),
    .Y(_0468_));
 sky130_fd_sc_hd__and4_1 _4348_ (.A(_0425_),
    .B(_1092_),
    .C(_1257_),
    .D(\A[1][4] ),
    .X(_0469_));
 sky130_fd_sc_hd__o21bai_1 _4349_ (.A1(_0467_),
    .A2(_0468_),
    .B1_N(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__nand3_1 _4350_ (.A(_0465_),
    .B(_0466_),
    .C(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__buf_2 _4351_ (.A(_0436_),
    .X(_0472_));
 sky130_fd_sc_hd__a22oi_1 _4352_ (.A1(_1312_),
    .A2(_0419_),
    .B1(_0472_),
    .B2(_1334_),
    .Y(_0473_));
 sky130_fd_sc_hd__and4_1 _4353_ (.A(\B[3][5] ),
    .B(_0419_),
    .C(_0436_),
    .D(\B[3][4] ),
    .X(_0474_));
 sky130_fd_sc_hd__nor2_1 _4354_ (.A(_0473_),
    .B(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__buf_2 _4355_ (.A(\A[1][1] ),
    .X(_0476_));
 sky130_fd_sc_hd__nand2_1 _4356_ (.A(_1587_),
    .B(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__xnor2_1 _4357_ (.A(_0475_),
    .B(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__a21o_1 _4358_ (.A1(_0465_),
    .A2(_0466_),
    .B1(_0470_),
    .X(_0479_));
 sky130_fd_sc_hd__nand3_1 _4359_ (.A(_0471_),
    .B(_0478_),
    .C(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__a21oi_1 _4360_ (.A1(_0442_),
    .A2(_0463_),
    .B1(_0462_),
    .Y(_0481_));
 sky130_fd_sc_hd__a211oi_1 _4361_ (.A1(_0471_),
    .A2(_0480_),
    .B1(_0464_),
    .C1(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__o21ba_1 _4362_ (.A1(_0437_),
    .A2(_0440_),
    .B1_N(_0438_),
    .X(_0483_));
 sky130_fd_sc_hd__o21ba_1 _4363_ (.A1(_0464_),
    .A2(_0482_),
    .B1_N(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__or3b_1 _4364_ (.A(_0464_),
    .B(_0482_),
    .C_N(_0483_),
    .X(_0485_));
 sky130_fd_sc_hd__and2b_1 _4365_ (.A_N(_0484_),
    .B(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__a31o_1 _4366_ (.A1(_0696_),
    .A2(_0421_),
    .A3(_0486_),
    .B1(_0484_),
    .X(_0487_));
 sky130_fd_sc_hd__nand2_1 _4367_ (.A(_0448_),
    .B(_0450_),
    .Y(_0488_));
 sky130_fd_sc_hd__clkbuf_4 _4368_ (.A(_0447_),
    .X(_0489_));
 sky130_fd_sc_hd__clkbuf_4 _4369_ (.A(_0454_),
    .X(_0490_));
 sky130_fd_sc_hd__a22o_1 _4370_ (.A1(_1959_),
    .A2(_0489_),
    .B1(_0490_),
    .B2(_0729_),
    .X(_0491_));
 sky130_fd_sc_hd__nand4_1 _4371_ (.A(_0740_),
    .B(_1959_),
    .C(_0489_),
    .D(_0490_),
    .Y(_0492_));
 sky130_fd_sc_hd__buf_2 _4372_ (.A(\A[0][4] ),
    .X(_0493_));
 sky130_fd_sc_hd__and4_1 _4373_ (.A(_0457_),
    .B(\B[1][3] ),
    .C(_0493_),
    .D(\B[1][4] ),
    .X(_0494_));
 sky130_fd_sc_hd__a22oi_1 _4374_ (.A1(_0927_),
    .A2(_0493_),
    .B1(_1026_),
    .B2(_0457_),
    .Y(_0495_));
 sky130_fd_sc_hd__and4bb_1 _4375_ (.A_N(_0494_),
    .B_N(_0495_),
    .C(\B[1][5] ),
    .D(_0455_),
    .X(_0496_));
 sky130_fd_sc_hd__a211o_1 _4376_ (.A1(_0491_),
    .A2(_0492_),
    .B1(_0494_),
    .C1(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__o211a_1 _4377_ (.A1(_0494_),
    .A2(_0496_),
    .B1(_0491_),
    .C1(_0492_),
    .X(_0498_));
 sky130_fd_sc_hd__a21oi_2 _4378_ (.A1(_0488_),
    .A2(_0497_),
    .B1(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__clkbuf_4 _4379_ (.A(_0430_),
    .X(_0500_));
 sky130_fd_sc_hd__nand2_1 _4380_ (.A(_1521_),
    .B(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__buf_2 _4381_ (.A(_0425_),
    .X(_0502_));
 sky130_fd_sc_hd__nand2_1 _4382_ (.A(_0502_),
    .B(_1543_),
    .Y(_0503_));
 sky130_fd_sc_hd__and4_1 _4383_ (.A(_0425_),
    .B(_1312_),
    .C(_0430_),
    .D(_1334_),
    .X(_0504_));
 sky130_fd_sc_hd__a21oi_1 _4384_ (.A1(_0501_),
    .A2(_0503_),
    .B1(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__clkbuf_4 _4385_ (.A(_0472_),
    .X(_0506_));
 sky130_fd_sc_hd__nand2_1 _4386_ (.A(_1587_),
    .B(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__xnor2_1 _4387_ (.A(_0505_),
    .B(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__nand2_1 _4388_ (.A(_0443_),
    .B(_1806_),
    .Y(_0509_));
 sky130_fd_sc_hd__nand2_1 _4389_ (.A(_0446_),
    .B(_2347_),
    .Y(_0510_));
 sky130_fd_sc_hd__a22o_1 _4390_ (.A1(\A[1][7] ),
    .A2(_1806_),
    .B1(_1202_),
    .B2(_0443_),
    .X(_0511_));
 sky130_fd_sc_hd__o21a_1 _4391_ (.A1(_0509_),
    .A2(_0510_),
    .B1(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__a21boi_2 _4392_ (.A1(_0424_),
    .A2(_0426_),
    .B1_N(_0423_),
    .Y(_0513_));
 sky130_fd_sc_hd__xnor2_1 _4393_ (.A(_0512_),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__xnor2_1 _4394_ (.A(_0508_),
    .B(_0514_),
    .Y(_0515_));
 sky130_fd_sc_hd__nor2_1 _4395_ (.A(_0499_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__nor3b_1 _4396_ (.A(_0434_),
    .B(_0435_),
    .C_N(_0441_),
    .Y(_0517_));
 sky130_fd_sc_hd__xor2_1 _4397_ (.A(_0499_),
    .B(_0515_),
    .X(_0518_));
 sky130_fd_sc_hd__o21a_1 _4398_ (.A1(_0434_),
    .A2(_0517_),
    .B1(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__a31oi_1 _4399_ (.A1(_2833_),
    .A2(_0506_),
    .A3(_0505_),
    .B1(_0504_),
    .Y(_0520_));
 sky130_fd_sc_hd__o21ba_1 _4400_ (.A1(_0516_),
    .A2(_0519_),
    .B1_N(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__or3b_1 _4401_ (.A(_0516_),
    .B(_0519_),
    .C_N(_0520_),
    .X(_0522_));
 sky130_fd_sc_hd__and2b_1 _4402_ (.A_N(_0521_),
    .B(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__nand2_1 _4403_ (.A(_0674_),
    .B(_0506_),
    .Y(_0524_));
 sky130_fd_sc_hd__xnor2_2 _4404_ (.A(_0523_),
    .B(_0524_),
    .Y(_0525_));
 sky130_fd_sc_hd__inv_2 _4405_ (.A(_0511_),
    .Y(_0526_));
 sky130_fd_sc_hd__nor2_1 _4406_ (.A(_0509_),
    .B(_0510_),
    .Y(_0527_));
 sky130_fd_sc_hd__nand2_1 _4407_ (.A(_0508_),
    .B(_0514_),
    .Y(_0528_));
 sky130_fd_sc_hd__o31ai_4 _4408_ (.A1(_0526_),
    .A2(_0527_),
    .A3(_0513_),
    .B1(_0528_),
    .Y(_0529_));
 sky130_fd_sc_hd__clkbuf_4 _4409_ (.A(_0740_),
    .X(_0530_));
 sky130_fd_sc_hd__clkbuf_4 _4410_ (.A(_0489_),
    .X(_0531_));
 sky130_fd_sc_hd__and4_1 _4411_ (.A(_0530_),
    .B(_2862_),
    .C(_0531_),
    .D(_0490_),
    .X(_0532_));
 sky130_fd_sc_hd__clkbuf_4 _4412_ (.A(_0457_),
    .X(_0533_));
 sky130_fd_sc_hd__a22oi_1 _4413_ (.A1(_1959_),
    .A2(_0490_),
    .B1(_0533_),
    .B2(_0729_),
    .Y(_0534_));
 sky130_fd_sc_hd__and4_1 _4414_ (.A(\B[1][6] ),
    .B(\B[1][7] ),
    .C(_0455_),
    .D(_0453_),
    .X(_0535_));
 sky130_fd_sc_hd__or2_1 _4415_ (.A(_0534_),
    .B(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__a22o_1 _4416_ (.A1(\A[0][5] ),
    .A2(_1015_),
    .B1(_0493_),
    .B2(_0938_),
    .X(_0537_));
 sky130_fd_sc_hd__and4_1 _4417_ (.A(\A[0][5] ),
    .B(\B[1][3] ),
    .C(_0493_),
    .D(_0938_),
    .X(_0538_));
 sky130_fd_sc_hd__a31o_1 _4418_ (.A1(_1904_),
    .A2(_0533_),
    .A3(_0537_),
    .B1(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__and2b_1 _4419_ (.A_N(_0536_),
    .B(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__and2b_1 _4420_ (.A_N(_0539_),
    .B(_0536_),
    .X(_0541_));
 sky130_fd_sc_hd__nor2_1 _4421_ (.A(_0540_),
    .B(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__a21o_1 _4422_ (.A1(_0532_),
    .A2(_0542_),
    .B1(_0540_),
    .X(_0543_));
 sky130_fd_sc_hd__and2_1 _4423_ (.A(_0443_),
    .B(_1312_),
    .X(_0544_));
 sky130_fd_sc_hd__inv_2 _4424_ (.A(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__clkbuf_4 _4425_ (.A(_0443_),
    .X(_0546_));
 sky130_fd_sc_hd__a22o_1 _4426_ (.A1(_0502_),
    .A2(_1521_),
    .B1(_1543_),
    .B2(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__o21a_1 _4427_ (.A1(_0503_),
    .A2(_0545_),
    .B1(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__nand2_1 _4428_ (.A(_1587_),
    .B(_0500_),
    .Y(_0549_));
 sky130_fd_sc_hd__xnor2_1 _4429_ (.A(_0548_),
    .B(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__and3_1 _4430_ (.A(_0446_),
    .B(_2347_),
    .C(_0509_),
    .X(_0551_));
 sky130_fd_sc_hd__xnor2_1 _4431_ (.A(_0550_),
    .B(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__xnor2_1 _4432_ (.A(_0543_),
    .B(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__xnor2_2 _4433_ (.A(_0529_),
    .B(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__buf_2 _4434_ (.A(\A[0][6] ),
    .X(_0555_));
 sky130_fd_sc_hd__buf_2 _4435_ (.A(\A[0][5] ),
    .X(_0556_));
 sky130_fd_sc_hd__a22o_1 _4436_ (.A1(_0555_),
    .A2(_0927_),
    .B1(_1026_),
    .B2(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__nand4_1 _4437_ (.A(_0555_),
    .B(_0556_),
    .C(_0927_),
    .D(_1026_),
    .Y(_0558_));
 sky130_fd_sc_hd__clkbuf_4 _4438_ (.A(net46),
    .X(_0559_));
 sky130_fd_sc_hd__and2_1 _4439_ (.A(\B[1][5] ),
    .B(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__a21o_1 _4440_ (.A1(_0557_),
    .A2(_0558_),
    .B1(_0560_),
    .X(_0561_));
 sky130_fd_sc_hd__nand3_1 _4441_ (.A(_0557_),
    .B(_0558_),
    .C(_0560_),
    .Y(_0562_));
 sky130_fd_sc_hd__nand2_1 _4442_ (.A(_0555_),
    .B(_2433_),
    .Y(_0563_));
 sky130_fd_sc_hd__and3_1 _4443_ (.A(\A[0][7] ),
    .B(_2432_),
    .C(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__and3_1 _4444_ (.A(_0561_),
    .B(_0562_),
    .C(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__and4_1 _4445_ (.A(\A[0][7] ),
    .B(\A[0][6] ),
    .C(_2496_),
    .D(\B[1][2] ),
    .X(_0566_));
 sky130_fd_sc_hd__clkbuf_4 _4446_ (.A(\A[0][7] ),
    .X(_0567_));
 sky130_fd_sc_hd__clkbuf_4 _4447_ (.A(net56),
    .X(_0568_));
 sky130_fd_sc_hd__and3_1 _4448_ (.A(_0567_),
    .B(_0568_),
    .C(_0949_),
    .X(_0569_));
 sky130_fd_sc_hd__a22o_1 _4449_ (.A1(_0567_),
    .A2(_2440_),
    .B1(_0949_),
    .B2(_0568_),
    .X(_0570_));
 sky130_fd_sc_hd__a21bo_1 _4450_ (.A1(_2440_),
    .A2(_0569_),
    .B1_N(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__clkbuf_4 _4451_ (.A(\A[0][5] ),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_4 _4452_ (.A(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__nand2_1 _4453_ (.A(_0573_),
    .B(_2856_),
    .Y(_0574_));
 sky130_fd_sc_hd__xor2_1 _4454_ (.A(_0571_),
    .B(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__o21ai_1 _4455_ (.A1(_0565_),
    .A2(_0566_),
    .B1(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__or3_1 _4456_ (.A(_0575_),
    .B(_0565_),
    .C(_0566_),
    .X(_0577_));
 sky130_fd_sc_hd__nand2_1 _4457_ (.A(_0576_),
    .B(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__a21bo_1 _4458_ (.A1(_0557_),
    .A2(_0560_),
    .B1_N(_0558_),
    .X(_0579_));
 sky130_fd_sc_hd__nand2_1 _4459_ (.A(_1959_),
    .B(_0533_),
    .Y(_0580_));
 sky130_fd_sc_hd__clkbuf_4 _4460_ (.A(_0559_),
    .X(_0581_));
 sky130_fd_sc_hd__nand2_1 _4461_ (.A(_0740_),
    .B(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__and4_1 _4462_ (.A(_0729_),
    .B(_1959_),
    .C(_0453_),
    .D(_0559_),
    .X(_0583_));
 sky130_fd_sc_hd__a21o_1 _4463_ (.A1(_0580_),
    .A2(_0582_),
    .B1(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__xnor2_1 _4464_ (.A(_0579_),
    .B(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__nor2_1 _4465_ (.A(_0535_),
    .B(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__and2_1 _4466_ (.A(_0535_),
    .B(_0585_),
    .X(_0587_));
 sky130_fd_sc_hd__or2_1 _4467_ (.A(_0586_),
    .B(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__xnor2_2 _4468_ (.A(_0578_),
    .B(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__a21oi_1 _4469_ (.A1(_0561_),
    .A2(_0562_),
    .B1(_0564_),
    .Y(_0590_));
 sky130_fd_sc_hd__and2b_1 _4470_ (.A_N(_0538_),
    .B(_0537_),
    .X(_0591_));
 sky130_fd_sc_hd__nand2_1 _4471_ (.A(_1904_),
    .B(_0533_),
    .Y(_0592_));
 sky130_fd_sc_hd__xnor2_2 _4472_ (.A(_0591_),
    .B(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__a22oi_1 _4473_ (.A1(\A[0][7] ),
    .A2(_2437_),
    .B1(_2438_),
    .B2(_0555_),
    .Y(_0594_));
 sky130_fd_sc_hd__or2_1 _4474_ (.A(_0566_),
    .B(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__and2_1 _4475_ (.A(_0556_),
    .B(_2438_),
    .X(_0596_));
 sky130_fd_sc_hd__a22o_1 _4476_ (.A1(\A[0][7] ),
    .A2(_2468_),
    .B1(_2437_),
    .B2(\A[0][6] ),
    .X(_0597_));
 sky130_fd_sc_hd__nand4_1 _4477_ (.A(\A[0][7] ),
    .B(_0555_),
    .C(_2468_),
    .D(_2437_),
    .Y(_0598_));
 sky130_fd_sc_hd__a21bo_1 _4478_ (.A1(_0596_),
    .A2(_0597_),
    .B1_N(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__xnor2_1 _4479_ (.A(_0595_),
    .B(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__or2b_1 _4480_ (.A(_0595_),
    .B_N(_0599_),
    .X(_0601_));
 sky130_fd_sc_hd__a21boi_1 _4481_ (.A1(_0593_),
    .A2(_0600_),
    .B1_N(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__xnor2_2 _4482_ (.A(_0532_),
    .B(_0542_),
    .Y(_0603_));
 sky130_fd_sc_hd__or2_1 _4483_ (.A(_0565_),
    .B(_0590_),
    .X(_0604_));
 sky130_fd_sc_hd__xnor2_1 _4484_ (.A(_0604_),
    .B(_0602_),
    .Y(_0605_));
 sky130_fd_sc_hd__o32a_1 _4485_ (.A1(_0565_),
    .A2(_0590_),
    .A3(_0602_),
    .B1(_0603_),
    .B2(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__xnor2_2 _4486_ (.A(_0589_),
    .B(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__xnor2_2 _4487_ (.A(_0554_),
    .B(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__nor3_1 _4488_ (.A(_0434_),
    .B(_0517_),
    .C(_0518_),
    .Y(_0609_));
 sky130_fd_sc_hd__nor2_1 _4489_ (.A(_0519_),
    .B(_0609_),
    .Y(_0610_));
 sky130_fd_sc_hd__xor2_2 _4490_ (.A(_0603_),
    .B(_0605_),
    .X(_0611_));
 sky130_fd_sc_hd__and2b_1 _4491_ (.A_N(_0498_),
    .B(_0497_),
    .X(_0612_));
 sky130_fd_sc_hd__xnor2_2 _4492_ (.A(_0488_),
    .B(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__xnor2_2 _4493_ (.A(_0593_),
    .B(_0600_),
    .Y(_0614_));
 sky130_fd_sc_hd__o2bb2a_1 _4494_ (.A1_N(_1904_),
    .A2_N(_0490_),
    .B1(_0494_),
    .B2(_0495_),
    .X(_0615_));
 sky130_fd_sc_hd__nor2_1 _4495_ (.A(_0496_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__nand3_1 _4496_ (.A(_0598_),
    .B(_0596_),
    .C(_0597_),
    .Y(_0617_));
 sky130_fd_sc_hd__a22o_1 _4497_ (.A1(_0572_),
    .A2(_2432_),
    .B1(_0598_),
    .B2(_0597_),
    .X(_0618_));
 sky130_fd_sc_hd__nand2_1 _4498_ (.A(_2438_),
    .B(_0493_),
    .Y(_0619_));
 sky130_fd_sc_hd__a22oi_2 _4499_ (.A1(\A[0][6] ),
    .A2(_2468_),
    .B1(_2437_),
    .B2(_0556_),
    .Y(_0620_));
 sky130_fd_sc_hd__and4_1 _4500_ (.A(\A[0][6] ),
    .B(\A[0][5] ),
    .C(_2470_),
    .D(_2496_),
    .X(_0621_));
 sky130_fd_sc_hd__o21bai_1 _4501_ (.A1(_0619_),
    .A2(_0620_),
    .B1_N(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__a21o_1 _4502_ (.A1(_0617_),
    .A2(_0618_),
    .B1(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__nand3_1 _4503_ (.A(_0617_),
    .B(_0618_),
    .C(_0622_),
    .Y(_0624_));
 sky130_fd_sc_hd__a21bo_1 _4504_ (.A1(_0616_),
    .A2(_0623_),
    .B1_N(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__xor2_2 _4505_ (.A(_0614_),
    .B(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__or2b_1 _4506_ (.A(_0614_),
    .B_N(_0625_),
    .X(_0627_));
 sky130_fd_sc_hd__o21a_1 _4507_ (.A1(_0613_),
    .A2(_0626_),
    .B1(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__xnor2_2 _4508_ (.A(_0611_),
    .B(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__or2b_1 _4509_ (.A(_0628_),
    .B_N(_0611_),
    .X(_0630_));
 sky130_fd_sc_hd__a21boi_2 _4510_ (.A1(_0610_),
    .A2(_0629_),
    .B1_N(_0630_),
    .Y(_0631_));
 sky130_fd_sc_hd__xor2_2 _4511_ (.A(_0608_),
    .B(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__xnor2_2 _4512_ (.A(_0525_),
    .B(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__nand2_1 _4513_ (.A(\B[3][7] ),
    .B(_0421_),
    .Y(_0634_));
 sky130_fd_sc_hd__xnor2_1 _4514_ (.A(_0486_),
    .B(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__xnor2_2 _4515_ (.A(_0610_),
    .B(_0629_),
    .Y(_0636_));
 sky130_fd_sc_hd__o211a_1 _4516_ (.A1(_0464_),
    .A2(_0481_),
    .B1(_0471_),
    .C1(_0480_),
    .X(_0637_));
 sky130_fd_sc_hd__nor2_1 _4517_ (.A(_0482_),
    .B(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__xnor2_2 _4518_ (.A(_0613_),
    .B(_0626_),
    .Y(_0639_));
 sky130_fd_sc_hd__and3_1 _4519_ (.A(_0445_),
    .B(_0461_),
    .C(_0460_),
    .X(_0640_));
 sky130_fd_sc_hd__a21oi_1 _4520_ (.A1(_0461_),
    .A2(_0460_),
    .B1(_0445_),
    .Y(_0641_));
 sky130_fd_sc_hd__or2_1 _4521_ (.A(_0640_),
    .B(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__nand3_1 _4522_ (.A(_0624_),
    .B(_0616_),
    .C(_0623_),
    .Y(_0643_));
 sky130_fd_sc_hd__a21o_1 _4523_ (.A1(_0624_),
    .A2(_0623_),
    .B1(_0616_),
    .X(_0644_));
 sky130_fd_sc_hd__nor2_1 _4524_ (.A(_0458_),
    .B(_0456_),
    .Y(_0645_));
 sky130_fd_sc_hd__xnor2_1 _4525_ (.A(_0452_),
    .B(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__or3_1 _4526_ (.A(_0621_),
    .B(_0619_),
    .C(_0620_),
    .X(_0647_));
 sky130_fd_sc_hd__o21ai_1 _4527_ (.A1(_0621_),
    .A2(_0620_),
    .B1(_0619_),
    .Y(_0648_));
 sky130_fd_sc_hd__nand2_1 _4528_ (.A(_2432_),
    .B(_0453_),
    .Y(_0649_));
 sky130_fd_sc_hd__a22oi_2 _4529_ (.A1(_0556_),
    .A2(_2468_),
    .B1(_2433_),
    .B2(_0559_),
    .Y(_0650_));
 sky130_fd_sc_hd__and4_1 _4530_ (.A(\A[0][5] ),
    .B(_2468_),
    .C(_2437_),
    .D(_0493_),
    .X(_0651_));
 sky130_fd_sc_hd__o21bai_1 _4531_ (.A1(_0649_),
    .A2(_0650_),
    .B1_N(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__a21o_1 _4532_ (.A1(_0647_),
    .A2(_0648_),
    .B1(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__nand3_1 _4533_ (.A(_0647_),
    .B(_0648_),
    .C(_0652_),
    .Y(_0654_));
 sky130_fd_sc_hd__a21bo_1 _4534_ (.A1(_0646_),
    .A2(_0653_),
    .B1_N(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__a21oi_1 _4535_ (.A1(_0643_),
    .A2(_0644_),
    .B1(_0655_),
    .Y(_0656_));
 sky130_fd_sc_hd__and3_1 _4536_ (.A(_0643_),
    .B(_0644_),
    .C(_0655_),
    .X(_0657_));
 sky130_fd_sc_hd__o21ba_1 _4537_ (.A1(_0642_),
    .A2(_0656_),
    .B1_N(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__xor2_2 _4538_ (.A(_0639_),
    .B(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__nor2_1 _4539_ (.A(_0639_),
    .B(_0658_),
    .Y(_0660_));
 sky130_fd_sc_hd__a21o_1 _4540_ (.A1(_0638_),
    .A2(_0659_),
    .B1(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__xnor2_1 _4541_ (.A(_0636_),
    .B(_0661_),
    .Y(_0662_));
 sky130_fd_sc_hd__or2b_1 _4542_ (.A(_0636_),
    .B_N(_0661_),
    .X(_0663_));
 sky130_fd_sc_hd__a21bo_1 _4543_ (.A1(_0635_),
    .A2(_0662_),
    .B1_N(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__xnor2_1 _4544_ (.A(_0633_),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__and2b_1 _4545_ (.A_N(_0633_),
    .B(_0664_),
    .X(_0666_));
 sky130_fd_sc_hd__a21o_1 _4546_ (.A1(_0487_),
    .A2(_0665_),
    .B1(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__a31oi_2 _4547_ (.A1(_0696_),
    .A2(_0506_),
    .A3(_0523_),
    .B1(_0521_),
    .Y(_0668_));
 sky130_fd_sc_hd__nor2_1 _4548_ (.A(_0608_),
    .B(_0631_),
    .Y(_0669_));
 sky130_fd_sc_hd__a21oi_1 _4549_ (.A1(_0525_),
    .A2(_0632_),
    .B1(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__buf_4 _4550_ (.A(_0500_),
    .X(_0671_));
 sky130_fd_sc_hd__nand2_1 _4551_ (.A(_0674_),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__nor2_1 _4552_ (.A(_0503_),
    .B(_0545_),
    .Y(_0673_));
 sky130_fd_sc_hd__a31o_1 _4553_ (.A1(_2833_),
    .A2(_0671_),
    .A3(_0547_),
    .B1(_0673_),
    .X(_0675_));
 sky130_fd_sc_hd__and2b_1 _4554_ (.A_N(_0552_),
    .B(_0543_),
    .X(_0676_));
 sky130_fd_sc_hd__a21o_1 _4555_ (.A1(_0529_),
    .A2(_0553_),
    .B1(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__xor2_1 _4556_ (.A(_0675_),
    .B(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__xor2_1 _4557_ (.A(_0672_),
    .B(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__or2_1 _4558_ (.A(_0589_),
    .B(_0606_),
    .X(_0680_));
 sky130_fd_sc_hd__o21ai_1 _4559_ (.A1(_0554_),
    .A2(_0607_),
    .B1(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__a21oi_1 _4560_ (.A1(_0550_),
    .A2(_0551_),
    .B1(_0527_),
    .Y(_0682_));
 sky130_fd_sc_hd__and2b_1 _4561_ (.A_N(_0584_),
    .B(_0579_),
    .X(_0683_));
 sky130_fd_sc_hd__clkbuf_4 _4562_ (.A(_0502_),
    .X(_0684_));
 sky130_fd_sc_hd__nand2_1 _4563_ (.A(_0684_),
    .B(_2833_),
    .Y(_0686_));
 sky130_fd_sc_hd__a21oi_1 _4564_ (.A1(_0446_),
    .A2(_2630_),
    .B1(_0544_),
    .Y(_0687_));
 sky130_fd_sc_hd__and3_1 _4565_ (.A(_0446_),
    .B(_2630_),
    .C(_0544_),
    .X(_0688_));
 sky130_fd_sc_hd__nor2_1 _4566_ (.A(_0687_),
    .B(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__xnor2_1 _4567_ (.A(_0686_),
    .B(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__o21a_1 _4568_ (.A1(_0683_),
    .A2(_0587_),
    .B1(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__nor3_1 _4569_ (.A(_0683_),
    .B(_0587_),
    .C(_0690_),
    .Y(_0692_));
 sky130_fd_sc_hd__nor2_1 _4570_ (.A(_0691_),
    .B(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__xnor2_1 _4571_ (.A(_0682_),
    .B(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__o21a_1 _4572_ (.A1(_0578_),
    .A2(_0588_),
    .B1(_0576_),
    .X(_0695_));
 sky130_fd_sc_hd__clkbuf_4 _4573_ (.A(_0568_),
    .X(_0697_));
 sky130_fd_sc_hd__clkbuf_4 _4574_ (.A(_0567_),
    .X(_0698_));
 sky130_fd_sc_hd__a22o_1 _4575_ (.A1(_0697_),
    .A2(_2856_),
    .B1(_0949_),
    .B2(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__nand2_1 _4576_ (.A(_2856_),
    .B(_0569_),
    .Y(_0700_));
 sky130_fd_sc_hd__nand2_1 _4577_ (.A(_0699_),
    .B(_0700_),
    .Y(_0701_));
 sky130_fd_sc_hd__a22o_1 _4578_ (.A1(_0572_),
    .A2(_0740_),
    .B1(_2862_),
    .B2(_0581_),
    .X(_0702_));
 sky130_fd_sc_hd__nand2_1 _4579_ (.A(_0572_),
    .B(_1959_),
    .Y(_0703_));
 sky130_fd_sc_hd__or2_1 _4580_ (.A(_0582_),
    .B(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__nand2_1 _4581_ (.A(_0702_),
    .B(_0704_),
    .Y(_0705_));
 sky130_fd_sc_hd__a32o_1 _4582_ (.A1(_0573_),
    .A2(_2856_),
    .A3(_0570_),
    .B1(_0569_),
    .B2(_2440_),
    .X(_0706_));
 sky130_fd_sc_hd__xor2_1 _4583_ (.A(_0705_),
    .B(_0706_),
    .X(_0708_));
 sky130_fd_sc_hd__xnor2_1 _4584_ (.A(_0583_),
    .B(_0708_),
    .Y(_0709_));
 sky130_fd_sc_hd__xnor2_1 _4585_ (.A(_0701_),
    .B(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__xnor2_1 _4586_ (.A(_0695_),
    .B(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__xnor2_1 _4587_ (.A(_0694_),
    .B(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__xnor2_1 _4588_ (.A(_0681_),
    .B(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__xor2_1 _4589_ (.A(_0679_),
    .B(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__xor2_1 _4590_ (.A(_0670_),
    .B(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__xnor2_2 _4591_ (.A(_0668_),
    .B(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__xnor2_1 _4592_ (.A(_0667_),
    .B(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__buf_2 _4593_ (.A(_0476_),
    .X(_0719_));
 sky130_fd_sc_hd__clkbuf_4 _4594_ (.A(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__and4_1 _4595_ (.A(_0447_),
    .B(_0454_),
    .C(_1015_),
    .D(_0938_),
    .X(_0721_));
 sky130_fd_sc_hd__a22oi_1 _4596_ (.A1(_0455_),
    .A2(_0927_),
    .B1(_1026_),
    .B2(_0447_),
    .Y(_0722_));
 sky130_fd_sc_hd__or2_1 _4597_ (.A(_0722_),
    .B(_0721_),
    .X(_0723_));
 sky130_fd_sc_hd__nand2_1 _4598_ (.A(_1904_),
    .B(_0444_),
    .Y(_0724_));
 sky130_fd_sc_hd__nor2_1 _4599_ (.A(_0723_),
    .B(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__clkbuf_4 _4600_ (.A(_0444_),
    .X(_0726_));
 sky130_fd_sc_hd__a22oi_1 _4601_ (.A1(_0740_),
    .A2(_0726_),
    .B1(_0784_),
    .B2(_0443_),
    .Y(_0727_));
 sky130_fd_sc_hd__nor2_1 _4602_ (.A(_0445_),
    .B(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__o21a_2 _4603_ (.A1(_0721_),
    .A2(_0725_),
    .B1(_0728_),
    .X(_0730_));
 sky130_fd_sc_hd__a21o_1 _4604_ (.A1(_0471_),
    .A2(_0479_),
    .B1(_0478_),
    .X(_0731_));
 sky130_fd_sc_hd__and3_1 _4605_ (.A(_0480_),
    .B(_0730_),
    .C(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__or3_1 _4606_ (.A(_0469_),
    .B(_0467_),
    .C(_0468_),
    .X(_0733_));
 sky130_fd_sc_hd__o21ai_1 _4607_ (.A1(_0469_),
    .A2(_0467_),
    .B1(_0468_),
    .Y(_0734_));
 sky130_fd_sc_hd__nand2_1 _4608_ (.A(_0419_),
    .B(_1202_),
    .Y(_0735_));
 sky130_fd_sc_hd__a22oi_2 _4609_ (.A1(_1103_),
    .A2(_0436_),
    .B1(\A[1][4] ),
    .B2(_1136_),
    .Y(_0736_));
 sky130_fd_sc_hd__and4_1 _4610_ (.A(_1092_),
    .B(_1257_),
    .C(_0436_),
    .D(\A[1][4] ),
    .X(_0737_));
 sky130_fd_sc_hd__o21bai_1 _4611_ (.A1(_0735_),
    .A2(_0736_),
    .B1_N(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__nand3_1 _4612_ (.A(_0733_),
    .B(_0734_),
    .C(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__a22oi_1 _4613_ (.A1(_1312_),
    .A2(_0476_),
    .B1(_0419_),
    .B2(_1543_),
    .Y(_0741_));
 sky130_fd_sc_hd__and4_1 _4614_ (.A(\B[3][5] ),
    .B(\A[1][1] ),
    .C(_0419_),
    .D(_1334_),
    .X(_0742_));
 sky130_fd_sc_hd__nor2_1 _4615_ (.A(_0741_),
    .B(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__nand2_1 _4616_ (.A(_1587_),
    .B(\A[1][0] ),
    .Y(_0744_));
 sky130_fd_sc_hd__xnor2_1 _4617_ (.A(_0743_),
    .B(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__a21o_1 _4618_ (.A1(_0733_),
    .A2(_0734_),
    .B1(_0738_),
    .X(_0746_));
 sky130_fd_sc_hd__nand3_1 _4619_ (.A(_0739_),
    .B(_0745_),
    .C(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__nand2_1 _4620_ (.A(_0739_),
    .B(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__nand3_1 _4621_ (.A(_0480_),
    .B(_0730_),
    .C(_0731_),
    .Y(_0749_));
 sky130_fd_sc_hd__a21o_1 _4622_ (.A1(_0480_),
    .A2(_0731_),
    .B1(_0730_),
    .X(_0750_));
 sky130_fd_sc_hd__and3_1 _4623_ (.A(_0748_),
    .B(_0749_),
    .C(_0750_),
    .X(_0752_));
 sky130_fd_sc_hd__o21ba_1 _4624_ (.A1(_0473_),
    .A2(_0477_),
    .B1_N(_0474_),
    .X(_0753_));
 sky130_fd_sc_hd__o21ba_1 _4625_ (.A1(_0732_),
    .A2(_0752_),
    .B1_N(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__or3b_1 _4626_ (.A(_0732_),
    .B(_0752_),
    .C_N(_0753_),
    .X(_0755_));
 sky130_fd_sc_hd__and2b_1 _4627_ (.A_N(_0754_),
    .B(_0755_),
    .X(_0756_));
 sky130_fd_sc_hd__a31o_1 _4628_ (.A1(_0685_),
    .A2(_0720_),
    .A3(_0756_),
    .B1(_0754_),
    .X(_0757_));
 sky130_fd_sc_hd__xor2_1 _4629_ (.A(_0635_),
    .B(_0662_),
    .X(_0758_));
 sky130_fd_sc_hd__nand2_1 _4630_ (.A(\B[3][7] ),
    .B(_0720_),
    .Y(_0759_));
 sky130_fd_sc_hd__xor2_2 _4631_ (.A(_0756_),
    .B(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__xnor2_1 _4632_ (.A(_0638_),
    .B(_0659_),
    .Y(_0761_));
 sky130_fd_sc_hd__a21oi_1 _4633_ (.A1(_0749_),
    .A2(_0750_),
    .B1(_0748_),
    .Y(_0763_));
 sky130_fd_sc_hd__nor2_1 _4634_ (.A(_0752_),
    .B(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__or3_1 _4635_ (.A(_0657_),
    .B(_0642_),
    .C(_0656_),
    .X(_0765_));
 sky130_fd_sc_hd__o21ai_2 _4636_ (.A1(_0657_),
    .A2(_0656_),
    .B1(_0642_),
    .Y(_0766_));
 sky130_fd_sc_hd__nand3_1 _4637_ (.A(_0654_),
    .B(_0646_),
    .C(_0653_),
    .Y(_0767_));
 sky130_fd_sc_hd__a21o_1 _4638_ (.A1(_0654_),
    .A2(_0653_),
    .B1(_0646_),
    .X(_0768_));
 sky130_fd_sc_hd__xor2_1 _4639_ (.A(_0723_),
    .B(_0724_),
    .X(_0769_));
 sky130_fd_sc_hd__or3_1 _4640_ (.A(_0651_),
    .B(_0649_),
    .C(_0650_),
    .X(_0770_));
 sky130_fd_sc_hd__o21ai_1 _4641_ (.A1(_0651_),
    .A2(_0650_),
    .B1(_0649_),
    .Y(_0771_));
 sky130_fd_sc_hd__nand2_1 _4642_ (.A(_0454_),
    .B(_2438_),
    .Y(_0772_));
 sky130_fd_sc_hd__a22oi_2 _4643_ (.A1(_2437_),
    .A2(_0457_),
    .B1(_0493_),
    .B2(_2468_),
    .Y(_0774_));
 sky130_fd_sc_hd__and4_1 _4644_ (.A(_2470_),
    .B(_2496_),
    .C(_0457_),
    .D(_0493_),
    .X(_0775_));
 sky130_fd_sc_hd__o21bai_1 _4645_ (.A1(_0772_),
    .A2(_0774_),
    .B1_N(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__a21o_1 _4646_ (.A1(_0770_),
    .A2(_0771_),
    .B1(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__nand3_1 _4647_ (.A(_0770_),
    .B(_0771_),
    .C(_0776_),
    .Y(_0778_));
 sky130_fd_sc_hd__a21bo_1 _4648_ (.A1(_0769_),
    .A2(_0777_),
    .B1_N(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__and3_1 _4649_ (.A(_0767_),
    .B(_0768_),
    .C(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__nand3_1 _4650_ (.A(_0767_),
    .B(_0768_),
    .C(_0779_),
    .Y(_0781_));
 sky130_fd_sc_hd__nor3_1 _4651_ (.A(_0721_),
    .B(_0725_),
    .C(_0728_),
    .Y(_0782_));
 sky130_fd_sc_hd__nor2_1 _4652_ (.A(_0730_),
    .B(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__a21o_1 _4653_ (.A1(_0767_),
    .A2(_0768_),
    .B1(_0779_),
    .X(_0785_));
 sky130_fd_sc_hd__and3_1 _4654_ (.A(_0781_),
    .B(_0783_),
    .C(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__a211o_1 _4655_ (.A1(_0765_),
    .A2(_0766_),
    .B1(_0780_),
    .C1(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__o211ai_4 _4656_ (.A1(_0780_),
    .A2(_0786_),
    .B1(_0765_),
    .C1(_0766_),
    .Y(_0788_));
 sky130_fd_sc_hd__a21boi_1 _4657_ (.A1(_0764_),
    .A2(_0787_),
    .B1_N(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__xnor2_1 _4658_ (.A(_0761_),
    .B(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__nor2_1 _4659_ (.A(_0761_),
    .B(_0789_),
    .Y(_0791_));
 sky130_fd_sc_hd__o21ba_1 _4660_ (.A1(_0760_),
    .A2(_0790_),
    .B1_N(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__xnor2_1 _4661_ (.A(_0758_),
    .B(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__and2b_1 _4662_ (.A_N(_0792_),
    .B(_0758_),
    .X(_0794_));
 sky130_fd_sc_hd__a21o_1 _4663_ (.A1(_0757_),
    .A2(_0793_),
    .B1(_0794_),
    .X(_0796_));
 sky130_fd_sc_hd__xor2_2 _4664_ (.A(_0487_),
    .B(_0665_),
    .X(_0797_));
 sky130_fd_sc_hd__and4_1 _4665_ (.A(_1521_),
    .B(\A[1][0] ),
    .C(_0476_),
    .D(_1543_),
    .X(_0798_));
 sky130_fd_sc_hd__and4_1 _4666_ (.A(\A[1][1] ),
    .B(_1136_),
    .C(_0419_),
    .D(_1257_),
    .X(_0799_));
 sky130_fd_sc_hd__a22oi_1 _4667_ (.A1(_1235_),
    .A2(_0419_),
    .B1(_1806_),
    .B2(\A[1][1] ),
    .Y(_0800_));
 sky130_fd_sc_hd__and4bb_1 _4668_ (.A_N(_0799_),
    .B_N(_0800_),
    .C(\A[1][0] ),
    .D(_1202_),
    .X(_0801_));
 sky130_fd_sc_hd__nor2_1 _4669_ (.A(_0799_),
    .B(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__nand2_1 _4670_ (.A(_0476_),
    .B(_2347_),
    .Y(_0803_));
 sky130_fd_sc_hd__and4_1 _4671_ (.A(_1092_),
    .B(\A[1][2] ),
    .C(\B[3][2] ),
    .D(\A[1][3] ),
    .X(_0804_));
 sky130_fd_sc_hd__a22o_1 _4672_ (.A1(\A[1][2] ),
    .A2(_1257_),
    .B1(_0436_),
    .B2(_1092_),
    .X(_0805_));
 sky130_fd_sc_hd__and2b_1 _4673_ (.A_N(_0804_),
    .B(_0805_),
    .X(_0807_));
 sky130_fd_sc_hd__xnor2_1 _4674_ (.A(_0803_),
    .B(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__and2b_1 _4675_ (.A_N(_0802_),
    .B(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__buf_2 _4676_ (.A(\A[1][0] ),
    .X(_0810_));
 sky130_fd_sc_hd__xnor2_1 _4677_ (.A(_0808_),
    .B(_0802_),
    .Y(_0811_));
 sky130_fd_sc_hd__and3_1 _4678_ (.A(_0810_),
    .B(_2630_),
    .C(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__a22oi_1 _4679_ (.A1(_1521_),
    .A2(\A[1][0] ),
    .B1(_0476_),
    .B2(_1543_),
    .Y(_0813_));
 sky130_fd_sc_hd__or2_1 _4680_ (.A(_0798_),
    .B(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__or3_1 _4681_ (.A(_0737_),
    .B(_0735_),
    .C(_0736_),
    .X(_0815_));
 sky130_fd_sc_hd__o21ai_1 _4682_ (.A1(_0737_),
    .A2(_0736_),
    .B1(_0735_),
    .Y(_0816_));
 sky130_fd_sc_hd__a31o_1 _4683_ (.A1(_0476_),
    .A2(_2347_),
    .A3(_0805_),
    .B1(_0804_),
    .X(_0818_));
 sky130_fd_sc_hd__and3_1 _4684_ (.A(_0815_),
    .B(_0816_),
    .C(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__a21oi_1 _4685_ (.A1(_0815_),
    .A2(_0816_),
    .B1(_0818_),
    .Y(_0820_));
 sky130_fd_sc_hd__nor2_1 _4686_ (.A(_0819_),
    .B(_0820_),
    .Y(_0821_));
 sky130_fd_sc_hd__xnor2_1 _4687_ (.A(_0814_),
    .B(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__o21a_1 _4688_ (.A1(_0809_),
    .A2(_0812_),
    .B1(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__and2_1 _4689_ (.A(_0798_),
    .B(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__or3_1 _4690_ (.A(_0775_),
    .B(_0772_),
    .C(_0774_),
    .X(_0825_));
 sky130_fd_sc_hd__o21ai_1 _4691_ (.A1(_0775_),
    .A2(_0774_),
    .B1(_0772_),
    .Y(_0826_));
 sky130_fd_sc_hd__nand2_1 _4692_ (.A(\A[0][1] ),
    .B(\B[1][2] ),
    .Y(_0827_));
 sky130_fd_sc_hd__a22oi_1 _4693_ (.A1(_2496_),
    .A2(\A[0][2] ),
    .B1(_0457_),
    .B2(_2470_),
    .Y(_0829_));
 sky130_fd_sc_hd__and4_1 _4694_ (.A(\B[1][0] ),
    .B(\B[1][1] ),
    .C(\A[0][2] ),
    .D(\A[0][3] ),
    .X(_0830_));
 sky130_fd_sc_hd__o21bai_1 _4695_ (.A1(_0827_),
    .A2(_0829_),
    .B1_N(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__nand3_1 _4696_ (.A(_0825_),
    .B(_0826_),
    .C(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__and4_1 _4697_ (.A(_0444_),
    .B(_0489_),
    .C(_2440_),
    .D(_0949_),
    .X(_0833_));
 sky130_fd_sc_hd__a22oi_1 _4698_ (.A1(_0531_),
    .A2(_2440_),
    .B1(_0949_),
    .B2(_0444_),
    .Y(_0834_));
 sky130_fd_sc_hd__nor2_1 _4699_ (.A(_0833_),
    .B(_0834_),
    .Y(_0835_));
 sky130_fd_sc_hd__a21o_1 _4700_ (.A1(_0825_),
    .A2(_0826_),
    .B1(_0831_),
    .X(_0836_));
 sky130_fd_sc_hd__nand3_1 _4701_ (.A(_0832_),
    .B(_0835_),
    .C(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__a21o_1 _4702_ (.A1(_0832_),
    .A2(_0836_),
    .B1(_0835_),
    .X(_0838_));
 sky130_fd_sc_hd__nand2_1 _4703_ (.A(_0726_),
    .B(_2440_),
    .Y(_0840_));
 sky130_fd_sc_hd__or3_1 _4704_ (.A(_0830_),
    .B(_0827_),
    .C(_0829_),
    .X(_0841_));
 sky130_fd_sc_hd__o21ai_1 _4705_ (.A1(_0830_),
    .A2(_0829_),
    .B1(_0827_),
    .Y(_0842_));
 sky130_fd_sc_hd__a22o_1 _4706_ (.A1(\A[0][1] ),
    .A2(_2496_),
    .B1(_0454_),
    .B2(_2470_),
    .X(_0843_));
 sky130_fd_sc_hd__and4_1 _4707_ (.A(_2470_),
    .B(\A[0][1] ),
    .C(\B[1][1] ),
    .D(\A[0][2] ),
    .X(_0844_));
 sky130_fd_sc_hd__a31o_1 _4708_ (.A1(\A[0][0] ),
    .A2(_2432_),
    .A3(_0843_),
    .B1(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__a21oi_2 _4709_ (.A1(_0841_),
    .A2(_0842_),
    .B1(_0845_),
    .Y(_0846_));
 sky130_fd_sc_hd__and3_1 _4710_ (.A(_0841_),
    .B(_0842_),
    .C(_0845_),
    .X(_0847_));
 sky130_fd_sc_hd__o21bai_2 _4711_ (.A1(_0840_),
    .A2(_0846_),
    .B1_N(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__nand3_4 _4712_ (.A(_0837_),
    .B(_0838_),
    .C(_0848_),
    .Y(_0849_));
 sky130_fd_sc_hd__a21o_1 _4713_ (.A1(_0837_),
    .A2(_0838_),
    .B1(_0848_),
    .X(_0851_));
 sky130_fd_sc_hd__nand4_4 _4714_ (.A(_2667_),
    .B(_0671_),
    .C(_0849_),
    .D(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__nand3_1 _4715_ (.A(_0778_),
    .B(_0769_),
    .C(_0777_),
    .Y(_0853_));
 sky130_fd_sc_hd__a21o_1 _4716_ (.A1(_0778_),
    .A2(_0777_),
    .B1(_0769_),
    .X(_0854_));
 sky130_fd_sc_hd__a21bo_1 _4717_ (.A1(_0835_),
    .A2(_0836_),
    .B1_N(_0832_),
    .X(_0855_));
 sky130_fd_sc_hd__and3_2 _4718_ (.A(_0853_),
    .B(_0854_),
    .C(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__and3_1 _4719_ (.A(_0502_),
    .B(_0784_),
    .C(_0833_),
    .X(_0857_));
 sky130_fd_sc_hd__a21oi_1 _4720_ (.A1(_0684_),
    .A2(_0784_),
    .B1(_0833_),
    .Y(_0858_));
 sky130_fd_sc_hd__or2_1 _4721_ (.A(_0857_),
    .B(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__a21oi_2 _4722_ (.A1(_0853_),
    .A2(_0854_),
    .B1(_0855_),
    .Y(_0860_));
 sky130_fd_sc_hd__nor3_4 _4723_ (.A(_0856_),
    .B(_0859_),
    .C(_0860_),
    .Y(_0862_));
 sky130_fd_sc_hd__o21a_1 _4724_ (.A1(_0856_),
    .A2(_0860_),
    .B1(_0859_),
    .X(_0863_));
 sky130_fd_sc_hd__a211oi_4 _4725_ (.A1(_0849_),
    .A2(_0852_),
    .B1(_0862_),
    .C1(_0863_),
    .Y(_0864_));
 sky130_fd_sc_hd__nor3_1 _4726_ (.A(_0822_),
    .B(_0809_),
    .C(_0812_),
    .Y(_0865_));
 sky130_fd_sc_hd__o211a_1 _4727_ (.A1(_0862_),
    .A2(_0863_),
    .B1(_0849_),
    .C1(_0852_),
    .X(_0866_));
 sky130_fd_sc_hd__nor4_2 _4728_ (.A(_0823_),
    .B(_0864_),
    .C(_0865_),
    .D(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__nand3_1 _4729_ (.A(_0781_),
    .B(_0783_),
    .C(_0785_),
    .Y(_0868_));
 sky130_fd_sc_hd__a21o_1 _4730_ (.A1(_0781_),
    .A2(_0785_),
    .B1(_0783_),
    .X(_0869_));
 sky130_fd_sc_hd__o211a_1 _4731_ (.A1(_0856_),
    .A2(_0862_),
    .B1(_0868_),
    .C1(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__o21ba_1 _4732_ (.A1(_0814_),
    .A2(_0820_),
    .B1_N(_0819_),
    .X(_0871_));
 sky130_fd_sc_hd__inv_2 _4733_ (.A(_0871_),
    .Y(_0873_));
 sky130_fd_sc_hd__a21o_1 _4734_ (.A1(_0739_),
    .A2(_0746_),
    .B1(_0745_),
    .X(_0874_));
 sky130_fd_sc_hd__nand3_1 _4735_ (.A(_0747_),
    .B(_0857_),
    .C(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__a21o_1 _4736_ (.A1(_0747_),
    .A2(_0874_),
    .B1(_0857_),
    .X(_0876_));
 sky130_fd_sc_hd__and3_1 _4737_ (.A(_0873_),
    .B(_0875_),
    .C(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__a21oi_1 _4738_ (.A1(_0875_),
    .A2(_0876_),
    .B1(_0873_),
    .Y(_0878_));
 sky130_fd_sc_hd__or2_1 _4739_ (.A(_0877_),
    .B(_0878_),
    .X(_0879_));
 sky130_fd_sc_hd__a211oi_2 _4740_ (.A1(_0868_),
    .A2(_0869_),
    .B1(_0856_),
    .C1(_0862_),
    .Y(_0880_));
 sky130_fd_sc_hd__or3_1 _4741_ (.A(_0870_),
    .B(_0879_),
    .C(_0880_),
    .X(_0881_));
 sky130_fd_sc_hd__o21ai_1 _4742_ (.A1(_0870_),
    .A2(_0880_),
    .B1(_0879_),
    .Y(_0882_));
 sky130_fd_sc_hd__o211a_1 _4743_ (.A1(_0864_),
    .A2(_0867_),
    .B1(_0881_),
    .C1(_0882_),
    .X(_0884_));
 sky130_fd_sc_hd__nor2_1 _4744_ (.A(_0798_),
    .B(_0823_),
    .Y(_0885_));
 sky130_fd_sc_hd__or2_1 _4745_ (.A(_0824_),
    .B(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__a211oi_1 _4746_ (.A1(_0881_),
    .A2(_0882_),
    .B1(_0864_),
    .C1(_0867_),
    .Y(_0887_));
 sky130_fd_sc_hd__nor3_2 _4747_ (.A(_0884_),
    .B(_0886_),
    .C(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__inv_2 _4748_ (.A(_0870_),
    .Y(_0889_));
 sky130_fd_sc_hd__and3_1 _4749_ (.A(_0788_),
    .B(_0764_),
    .C(_0787_),
    .X(_0890_));
 sky130_fd_sc_hd__a21oi_1 _4750_ (.A1(_0788_),
    .A2(_0787_),
    .B1(_0764_),
    .Y(_0891_));
 sky130_fd_sc_hd__a211oi_1 _4751_ (.A1(_0889_),
    .A2(_0881_),
    .B1(_0890_),
    .C1(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__and3_1 _4752_ (.A(_0747_),
    .B(_0857_),
    .C(_0874_),
    .X(_0893_));
 sky130_fd_sc_hd__o21ba_1 _4753_ (.A1(_0741_),
    .A2(_0744_),
    .B1_N(_0742_),
    .X(_0895_));
 sky130_fd_sc_hd__o21ba_1 _4754_ (.A1(_0893_),
    .A2(_0877_),
    .B1_N(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__or3b_1 _4755_ (.A(_0893_),
    .B(_0877_),
    .C_N(_0895_),
    .X(_0897_));
 sky130_fd_sc_hd__and2b_1 _4756_ (.A_N(_0896_),
    .B(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__clkbuf_4 _4757_ (.A(_0810_),
    .X(_0899_));
 sky130_fd_sc_hd__nand2_1 _4758_ (.A(_0674_),
    .B(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__xor2_1 _4759_ (.A(_0898_),
    .B(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__o211a_1 _4760_ (.A1(_0890_),
    .A2(_0891_),
    .B1(_0889_),
    .C1(_0881_),
    .X(_0902_));
 sky130_fd_sc_hd__or3_1 _4761_ (.A(_0892_),
    .B(_0901_),
    .C(_0902_),
    .X(_0903_));
 sky130_fd_sc_hd__o21ai_1 _4762_ (.A1(_0892_),
    .A2(_0902_),
    .B1(_0901_),
    .Y(_0904_));
 sky130_fd_sc_hd__o211ai_1 _4763_ (.A1(_0884_),
    .A2(_0888_),
    .B1(_0903_),
    .C1(_0904_),
    .Y(_0906_));
 sky130_fd_sc_hd__a211o_1 _4764_ (.A1(_0903_),
    .A2(_0904_),
    .B1(_0884_),
    .C1(_0888_),
    .X(_0907_));
 sky130_fd_sc_hd__nand3_1 _4765_ (.A(_0824_),
    .B(_0906_),
    .C(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__a21o_1 _4766_ (.A1(_0906_),
    .A2(_0907_),
    .B1(_0824_),
    .X(_0909_));
 sky130_fd_sc_hd__a22o_1 _4767_ (.A1(_2667_),
    .A2(_0671_),
    .B1(_0849_),
    .B2(_0851_),
    .X(_0910_));
 sky130_fd_sc_hd__and2_1 _4768_ (.A(_2667_),
    .B(_0506_),
    .X(_0911_));
 sky130_fd_sc_hd__or3_1 _4769_ (.A(_0840_),
    .B(_0847_),
    .C(_0846_),
    .X(_0912_));
 sky130_fd_sc_hd__o21ai_1 _4770_ (.A1(_0847_),
    .A2(_0846_),
    .B1(_0840_),
    .Y(_0913_));
 sky130_fd_sc_hd__nand2_1 _4771_ (.A(_0444_),
    .B(_2432_),
    .Y(_0914_));
 sky130_fd_sc_hd__and2b_1 _4772_ (.A_N(_0844_),
    .B(_0843_),
    .X(_0915_));
 sky130_fd_sc_hd__xnor2_1 _4773_ (.A(_0914_),
    .B(_0915_),
    .Y(_0917_));
 sky130_fd_sc_hd__and4_1 _4774_ (.A(_0726_),
    .B(_2471_),
    .C(_0531_),
    .D(_2433_),
    .X(_0918_));
 sky130_fd_sc_hd__and2_1 _4775_ (.A(_0917_),
    .B(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__a21o_1 _4776_ (.A1(_0912_),
    .A2(_0913_),
    .B1(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__nand3_1 _4777_ (.A(_0912_),
    .B(_0919_),
    .C(_0913_),
    .Y(_0921_));
 sky130_fd_sc_hd__a21bo_1 _4778_ (.A1(_0911_),
    .A2(_0920_),
    .B1_N(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__nand3_2 _4779_ (.A(_0852_),
    .B(_0910_),
    .C(_0922_),
    .Y(_0923_));
 sky130_fd_sc_hd__and3_1 _4780_ (.A(_0852_),
    .B(_0910_),
    .C(_0922_),
    .X(_0924_));
 sky130_fd_sc_hd__nand2_1 _4781_ (.A(_0810_),
    .B(_2630_),
    .Y(_0925_));
 sky130_fd_sc_hd__xnor2_1 _4782_ (.A(_0925_),
    .B(_0811_),
    .Y(_0926_));
 sky130_fd_sc_hd__o2bb2a_1 _4783_ (.A1_N(\A[1][0] ),
    .A2_N(_2347_),
    .B1(_0799_),
    .B2(_0800_),
    .X(_0928_));
 sky130_fd_sc_hd__nor2_1 _4784_ (.A(_0801_),
    .B(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__and4_1 _4785_ (.A(\A[1][0] ),
    .B(_0719_),
    .C(_1235_),
    .D(_1806_),
    .X(_0930_));
 sky130_fd_sc_hd__and2_1 _4786_ (.A(_0929_),
    .B(_0930_),
    .X(_0931_));
 sky130_fd_sc_hd__and2_1 _4787_ (.A(_0926_),
    .B(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__nor2_1 _4788_ (.A(_0926_),
    .B(_0931_),
    .Y(_0933_));
 sky130_fd_sc_hd__or2_1 _4789_ (.A(_0932_),
    .B(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__a21oi_1 _4790_ (.A1(_0852_),
    .A2(_0910_),
    .B1(_0922_),
    .Y(_0935_));
 sky130_fd_sc_hd__or3_1 _4791_ (.A(_0924_),
    .B(_0934_),
    .C(_0935_),
    .X(_0936_));
 sky130_fd_sc_hd__o22a_1 _4792_ (.A1(_0823_),
    .A2(_0865_),
    .B1(_0866_),
    .B2(_0864_),
    .X(_0937_));
 sky130_fd_sc_hd__a211o_1 _4793_ (.A1(_0923_),
    .A2(_0936_),
    .B1(_0867_),
    .C1(_0937_),
    .X(_0939_));
 sky130_fd_sc_hd__o211ai_2 _4794_ (.A1(_0867_),
    .A2(_0937_),
    .B1(_0923_),
    .C1(_0936_),
    .Y(_0940_));
 sky130_fd_sc_hd__nand3_2 _4795_ (.A(_0932_),
    .B(_0939_),
    .C(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__o21a_1 _4796_ (.A1(_0884_),
    .A2(_0887_),
    .B1(_0886_),
    .X(_0942_));
 sky130_fd_sc_hd__a211oi_2 _4797_ (.A1(_0939_),
    .A2(_0941_),
    .B1(_0942_),
    .C1(_0888_),
    .Y(_0943_));
 sky130_fd_sc_hd__a21oi_1 _4798_ (.A1(_0908_),
    .A2(_0909_),
    .B1(_0943_),
    .Y(_0944_));
 sky130_fd_sc_hd__o21ai_1 _4799_ (.A1(_0924_),
    .A2(_0935_),
    .B1(_0934_),
    .Y(_0945_));
 sky130_fd_sc_hd__nand3_1 _4800_ (.A(_0921_),
    .B(_0911_),
    .C(_0920_),
    .Y(_0946_));
 sky130_fd_sc_hd__a21o_1 _4801_ (.A1(_0921_),
    .A2(_0920_),
    .B1(_0911_),
    .X(_0947_));
 sky130_fd_sc_hd__xor2_1 _4802_ (.A(_0917_),
    .B(_0918_),
    .X(_0948_));
 sky130_fd_sc_hd__and3_1 _4803_ (.A(_2667_),
    .B(_0421_),
    .C(_0948_),
    .X(_0950_));
 sky130_fd_sc_hd__a21o_1 _4804_ (.A1(_0946_),
    .A2(_0947_),
    .B1(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__nor2_1 _4805_ (.A(_0929_),
    .B(_0930_),
    .Y(_0952_));
 sky130_fd_sc_hd__nor2_1 _4806_ (.A(_0931_),
    .B(_0952_),
    .Y(_0953_));
 sky130_fd_sc_hd__and3_1 _4807_ (.A(_0946_),
    .B(_0947_),
    .C(_0950_),
    .X(_0954_));
 sky130_fd_sc_hd__a21o_1 _4808_ (.A1(_0951_),
    .A2(_0953_),
    .B1(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__and3_1 _4809_ (.A(_0936_),
    .B(_0945_),
    .C(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__a21o_1 _4810_ (.A1(_0936_),
    .A2(_0945_),
    .B1(_0955_),
    .X(_0957_));
 sky130_fd_sc_hd__and2b_1 _4811_ (.A_N(_0956_),
    .B(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__or2b_1 _4812_ (.A(_0954_),
    .B_N(_0951_),
    .X(_0959_));
 sky130_fd_sc_hd__xnor2_2 _4813_ (.A(_0959_),
    .B(_0953_),
    .Y(_0961_));
 sky130_fd_sc_hd__a21oi_1 _4814_ (.A1(_2667_),
    .A2(_0421_),
    .B1(_0948_),
    .Y(_0962_));
 sky130_fd_sc_hd__nor2_1 _4815_ (.A(_0950_),
    .B(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__buf_4 _4816_ (.A(_0444_),
    .X(_0964_));
 sky130_fd_sc_hd__a22oi_1 _4817_ (.A1(_2471_),
    .A2(_0531_),
    .B1(_2433_),
    .B2(_0964_),
    .Y(_0965_));
 sky130_fd_sc_hd__nor2_1 _4818_ (.A(_0918_),
    .B(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__and3_1 _4819_ (.A(_2778_),
    .B(_0719_),
    .C(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__xnor2_1 _4820_ (.A(_0963_),
    .B(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__a22oi_1 _4821_ (.A1(_0720_),
    .A2(_1235_),
    .B1(_1806_),
    .B2(_0810_),
    .Y(_0969_));
 sky130_fd_sc_hd__or2_1 _4822_ (.A(_0930_),
    .B(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__or2_1 _4823_ (.A(_0968_),
    .B(_0970_),
    .X(_0972_));
 sky130_fd_sc_hd__a21bo_1 _4824_ (.A1(_0963_),
    .A2(_0967_),
    .B1_N(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__xor2_1 _4825_ (.A(_0961_),
    .B(_0973_),
    .X(_0974_));
 sky130_fd_sc_hd__nand2_1 _4826_ (.A(_0968_),
    .B(_0970_),
    .Y(_0975_));
 sky130_fd_sc_hd__a21oi_1 _4827_ (.A1(_2778_),
    .A2(_0720_),
    .B1(_0966_),
    .Y(_0976_));
 sky130_fd_sc_hd__nor2_1 _4828_ (.A(_0967_),
    .B(_0976_),
    .Y(_0977_));
 sky130_fd_sc_hd__and4_1 _4829_ (.A(_0964_),
    .B(_0810_),
    .C(_2471_),
    .D(_2778_),
    .X(_0978_));
 sky130_fd_sc_hd__nand2_1 _4830_ (.A(_0899_),
    .B(_1235_),
    .Y(_0979_));
 sky130_fd_sc_hd__xnor2_1 _4831_ (.A(_0977_),
    .B(_0978_),
    .Y(_0980_));
 sky130_fd_sc_hd__nor2_1 _4832_ (.A(_0979_),
    .B(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__a21o_1 _4833_ (.A1(_0977_),
    .A2(_0978_),
    .B1(_0981_),
    .X(_0983_));
 sky130_fd_sc_hd__and3_1 _4834_ (.A(_0972_),
    .B(_0975_),
    .C(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__nand3_1 _4835_ (.A(_0958_),
    .B(_0974_),
    .C(_0984_),
    .Y(_0985_));
 sky130_fd_sc_hd__a21o_1 _4836_ (.A1(_0939_),
    .A2(_0940_),
    .B1(_0932_),
    .X(_0986_));
 sky130_fd_sc_hd__a31o_1 _4837_ (.A1(_0957_),
    .A2(_0961_),
    .A3(_0973_),
    .B1(_0956_),
    .X(_0987_));
 sky130_fd_sc_hd__and3_1 _4838_ (.A(_0941_),
    .B(_0986_),
    .C(_0987_),
    .X(_0988_));
 sky130_fd_sc_hd__a21oi_1 _4839_ (.A1(_0941_),
    .A2(_0986_),
    .B1(_0987_),
    .Y(_0989_));
 sky130_fd_sc_hd__or3_1 _4840_ (.A(_0985_),
    .B(_0988_),
    .C(_0989_),
    .X(_0990_));
 sky130_fd_sc_hd__nand2_1 _4841_ (.A(_0961_),
    .B(_0973_),
    .Y(_0991_));
 sky130_fd_sc_hd__and2_1 _4842_ (.A(_0941_),
    .B(_0986_),
    .X(_0992_));
 sky130_fd_sc_hd__or4bb_1 _4843_ (.A(_0956_),
    .B(_0991_),
    .C_N(_0992_),
    .D_N(_0957_),
    .X(_0994_));
 sky130_fd_sc_hd__o211a_1 _4844_ (.A1(_0888_),
    .A2(_0942_),
    .B1(_0941_),
    .C1(_0939_),
    .X(_0995_));
 sky130_fd_sc_hd__and4bb_1 _4845_ (.A_N(_0943_),
    .B_N(_0995_),
    .C(_0992_),
    .D(_0956_),
    .X(_0996_));
 sky130_fd_sc_hd__o2bb2a_1 _4846_ (.A1_N(_0956_),
    .A2_N(_0992_),
    .B1(_0995_),
    .B2(_0943_),
    .X(_0997_));
 sky130_fd_sc_hd__a211o_1 _4847_ (.A1(_0990_),
    .A2(_0994_),
    .B1(_0996_),
    .C1(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__o211ai_1 _4848_ (.A1(_0943_),
    .A2(_0996_),
    .B1(_0908_),
    .C1(_0909_),
    .Y(_0999_));
 sky130_fd_sc_hd__o21a_1 _4849_ (.A1(_0944_),
    .A2(_0998_),
    .B1(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__xnor2_1 _4850_ (.A(_0757_),
    .B(_0793_),
    .Y(_1001_));
 sky130_fd_sc_hd__a31o_1 _4851_ (.A1(_0685_),
    .A2(_0899_),
    .A3(_0898_),
    .B1(_0896_),
    .X(_1002_));
 sky130_fd_sc_hd__xor2_2 _4852_ (.A(_0760_),
    .B(_0790_),
    .X(_1003_));
 sky130_fd_sc_hd__o21bai_2 _4853_ (.A1(_0901_),
    .A2(_0902_),
    .B1_N(_0892_),
    .Y(_1005_));
 sky130_fd_sc_hd__xor2_2 _4854_ (.A(_1003_),
    .B(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__and2_1 _4855_ (.A(_1003_),
    .B(_1005_),
    .X(_1007_));
 sky130_fd_sc_hd__a21oi_1 _4856_ (.A1(_1002_),
    .A2(_1006_),
    .B1(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__xnor2_1 _4857_ (.A(_1001_),
    .B(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__xor2_2 _4858_ (.A(_1002_),
    .B(_1006_),
    .X(_1010_));
 sky130_fd_sc_hd__a21boi_1 _4859_ (.A1(_0824_),
    .A2(_0907_),
    .B1_N(_0906_),
    .Y(_1011_));
 sky130_fd_sc_hd__xor2_2 _4860_ (.A(_1010_),
    .B(_1011_),
    .X(_1012_));
 sky130_fd_sc_hd__or2_1 _4861_ (.A(_1009_),
    .B(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__nor2_1 _4862_ (.A(_1000_),
    .B(_1013_),
    .Y(_1014_));
 sky130_fd_sc_hd__or2_1 _4863_ (.A(_1001_),
    .B(_1008_),
    .X(_1016_));
 sky130_fd_sc_hd__or2b_1 _4864_ (.A(_1011_),
    .B_N(_1010_),
    .X(_1017_));
 sky130_fd_sc_hd__and2_1 _4865_ (.A(_1001_),
    .B(_1008_),
    .X(_1018_));
 sky130_fd_sc_hd__a21oi_1 _4866_ (.A1(_1016_),
    .A2(_1017_),
    .B1(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__xor2_1 _4867_ (.A(_0796_),
    .B(_0797_),
    .X(_1020_));
 sky130_fd_sc_hd__o21ai_1 _4868_ (.A1(_1014_),
    .A2(_1019_),
    .B1(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__a21boi_1 _4869_ (.A1(_0796_),
    .A2(_0797_),
    .B1_N(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__xor2_1 _4870_ (.A(_0717_),
    .B(_1022_),
    .X(_1023_));
 sky130_fd_sc_hd__nor2_2 _4871_ (.A(net15),
    .B(_2883_),
    .Y(_1024_));
 sky130_fd_sc_hd__clkbuf_4 _4872_ (.A(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__a221o_1 _4873_ (.A1(_2885_),
    .A2(_0418_),
    .B1(_1023_),
    .B2(_2882_),
    .C1(_1025_),
    .X(_1027_));
 sky130_fd_sc_hd__clkbuf_4 _4874_ (.A(net1),
    .X(_1028_));
 sky130_fd_sc_hd__buf_4 _4875_ (.A(_0079_),
    .X(_1029_));
 sky130_fd_sc_hd__and3_1 _4876_ (.A(_2887_),
    .B(_2964_),
    .C(_0489_),
    .X(_1030_));
 sky130_fd_sc_hd__a22o_1 _4877_ (.A1(_2964_),
    .A2(_0444_),
    .B1(_0489_),
    .B2(_2887_),
    .X(_1031_));
 sky130_fd_sc_hd__a21bo_1 _4878_ (.A1(_0726_),
    .A2(_1030_),
    .B1_N(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__nand2_1 _4879_ (.A(_0446_),
    .B(_0085_),
    .Y(_1033_));
 sky130_fd_sc_hd__xnor2_1 _4880_ (.A(_1032_),
    .B(_1033_),
    .Y(_1034_));
 sky130_fd_sc_hd__and4_1 _4881_ (.A(_0455_),
    .B(_0453_),
    .C(_0152_),
    .D(_0153_),
    .X(_1035_));
 sky130_fd_sc_hd__a22oi_1 _4882_ (.A1(_0533_),
    .A2(_0152_),
    .B1(_0153_),
    .B2(_0490_),
    .Y(_1036_));
 sky130_fd_sc_hd__and4bb_1 _4883_ (.A_N(_1035_),
    .B_N(_1036_),
    .C(_2988_),
    .D(_0531_),
    .X(_1038_));
 sky130_fd_sc_hd__or2_1 _4884_ (.A(_1035_),
    .B(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__or2b_1 _4885_ (.A(_1034_),
    .B_N(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__xnor2_2 _4886_ (.A(_1039_),
    .B(_1034_),
    .Y(_1041_));
 sky130_fd_sc_hd__and4_1 _4887_ (.A(_2888_),
    .B(_0443_),
    .C(_0726_),
    .D(_0085_),
    .X(_1042_));
 sky130_fd_sc_hd__nand2_1 _4888_ (.A(_1041_),
    .B(_1042_),
    .Y(_1043_));
 sky130_fd_sc_hd__a22oi_1 _4889_ (.A1(_0159_),
    .A2(_0472_),
    .B1(_0500_),
    .B2(_0160_),
    .Y(_1044_));
 sky130_fd_sc_hd__and4_1 _4890_ (.A(_0159_),
    .B(_0472_),
    .C(_0500_),
    .D(_2917_),
    .X(_1045_));
 sky130_fd_sc_hd__nor2_1 _4891_ (.A(_1044_),
    .B(_1045_),
    .Y(_1046_));
 sky130_fd_sc_hd__nand2_1 _4892_ (.A(_2921_),
    .B(_0420_),
    .Y(_1047_));
 sky130_fd_sc_hd__xnor2_1 _4893_ (.A(_1046_),
    .B(_1047_),
    .Y(_1049_));
 sky130_fd_sc_hd__inv_2 _4894_ (.A(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__and3_1 _4895_ (.A(_0422_),
    .B(_0221_),
    .C(_0220_),
    .X(_1051_));
 sky130_fd_sc_hd__a22o_1 _4896_ (.A1(\A[1][7] ),
    .A2(_0221_),
    .B1(_0220_),
    .B2(_0422_),
    .X(_1052_));
 sky130_fd_sc_hd__a21bo_1 _4897_ (.A1(_0446_),
    .A2(_1051_),
    .B1_N(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__nand2_1 _4898_ (.A(_0502_),
    .B(_3002_),
    .Y(_1054_));
 sky130_fd_sc_hd__xor2_1 _4899_ (.A(_1053_),
    .B(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__a22o_1 _4900_ (.A1(_0422_),
    .A2(_0221_),
    .B1(_0220_),
    .B2(_0425_),
    .X(_1056_));
 sky130_fd_sc_hd__and4_1 _4901_ (.A(_0422_),
    .B(_0425_),
    .C(_2903_),
    .D(_2905_),
    .X(_1057_));
 sky130_fd_sc_hd__a31o_1 _4902_ (.A1(_3002_),
    .A2(_0500_),
    .A3(_1056_),
    .B1(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__xnor2_1 _4903_ (.A(_1055_),
    .B(_1058_),
    .Y(_1060_));
 sky130_fd_sc_hd__xnor2_1 _4904_ (.A(_1050_),
    .B(_1060_),
    .Y(_1061_));
 sky130_fd_sc_hd__a21oi_1 _4905_ (.A1(_1040_),
    .A2(_1043_),
    .B1(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__a22oi_1 _4906_ (.A1(_0378_),
    .A2(_0420_),
    .B1(_0472_),
    .B2(_0229_),
    .Y(_1063_));
 sky130_fd_sc_hd__and4_1 _4907_ (.A(_0159_),
    .B(_0420_),
    .C(_0472_),
    .D(_0160_),
    .X(_1064_));
 sky130_fd_sc_hd__nor2_1 _4908_ (.A(_1063_),
    .B(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__nand2_1 _4909_ (.A(_2921_),
    .B(_0719_),
    .Y(_1066_));
 sky130_fd_sc_hd__xnor2_1 _4910_ (.A(_1065_),
    .B(_1066_),
    .Y(_1067_));
 sky130_fd_sc_hd__and2b_1 _4911_ (.A_N(_1057_),
    .B(_1056_),
    .X(_1068_));
 sky130_fd_sc_hd__nand2_1 _4912_ (.A(_3002_),
    .B(_0500_),
    .Y(_1069_));
 sky130_fd_sc_hd__xnor2_1 _4913_ (.A(_1068_),
    .B(_1069_),
    .Y(_1071_));
 sky130_fd_sc_hd__and4_1 _4914_ (.A(_0425_),
    .B(_0221_),
    .C(_2905_),
    .D(_0430_),
    .X(_1072_));
 sky130_fd_sc_hd__a22oi_1 _4915_ (.A1(_0425_),
    .A2(_0221_),
    .B1(_0294_),
    .B2(_0430_),
    .Y(_1073_));
 sky130_fd_sc_hd__and4bb_1 _4916_ (.A_N(_1072_),
    .B_N(_1073_),
    .C(_0472_),
    .D(_3001_),
    .X(_1074_));
 sky130_fd_sc_hd__nor2_1 _4917_ (.A(_1072_),
    .B(_1074_),
    .Y(_1075_));
 sky130_fd_sc_hd__xnor2_1 _4918_ (.A(_1071_),
    .B(_1075_),
    .Y(_1076_));
 sky130_fd_sc_hd__and2b_1 _4919_ (.A_N(_1075_),
    .B(_1071_),
    .X(_1077_));
 sky130_fd_sc_hd__a21oi_1 _4920_ (.A1(_1067_),
    .A2(_1076_),
    .B1(_1077_),
    .Y(_1078_));
 sky130_fd_sc_hd__and3_1 _4921_ (.A(_1040_),
    .B(_1043_),
    .C(_1061_),
    .X(_1079_));
 sky130_fd_sc_hd__nor2_1 _4922_ (.A(_1062_),
    .B(_1079_),
    .Y(_1080_));
 sky130_fd_sc_hd__and2b_1 _4923_ (.A_N(_1078_),
    .B(_1080_),
    .X(_1082_));
 sky130_fd_sc_hd__o21ba_1 _4924_ (.A1(_1044_),
    .A2(_1047_),
    .B1_N(_1045_),
    .X(_1083_));
 sky130_fd_sc_hd__o21ba_1 _4925_ (.A1(_1062_),
    .A2(_1082_),
    .B1_N(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__or3b_1 _4926_ (.A(_1062_),
    .B(_1082_),
    .C_N(_1083_),
    .X(_1085_));
 sky130_fd_sc_hd__and2b_1 _4927_ (.A_N(_1084_),
    .B(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__a31o_1 _4928_ (.A1(_1029_),
    .A2(_0421_),
    .A3(_1086_),
    .B1(_1084_),
    .X(_1087_));
 sky130_fd_sc_hd__nand4_1 _4929_ (.A(_0567_),
    .B(_0568_),
    .C(_0280_),
    .D(_0282_),
    .Y(_1088_));
 sky130_fd_sc_hd__a22o_1 _4930_ (.A1(_0567_),
    .A2(_0279_),
    .B1(_0282_),
    .B2(_0568_),
    .X(_1089_));
 sky130_fd_sc_hd__and2_1 _4931_ (.A(_0572_),
    .B(_0241_),
    .X(_1090_));
 sky130_fd_sc_hd__nand3_1 _4932_ (.A(_1088_),
    .B(_1089_),
    .C(_1090_),
    .Y(_1091_));
 sky130_fd_sc_hd__a21o_1 _4933_ (.A1(_1088_),
    .A2(_1089_),
    .B1(_1090_),
    .X(_1093_));
 sky130_fd_sc_hd__a22oi_2 _4934_ (.A1(_0555_),
    .A2(_0279_),
    .B1(_0282_),
    .B2(_0572_),
    .Y(_1094_));
 sky130_fd_sc_hd__nand2_1 _4935_ (.A(_0241_),
    .B(_0581_),
    .Y(_1095_));
 sky130_fd_sc_hd__and4_1 _4936_ (.A(_0555_),
    .B(_0556_),
    .C(_0279_),
    .D(_0281_),
    .X(_1096_));
 sky130_fd_sc_hd__o21bai_1 _4937_ (.A1(_1094_),
    .A2(_1095_),
    .B1_N(_1096_),
    .Y(_1097_));
 sky130_fd_sc_hd__nand3_2 _4938_ (.A(_1091_),
    .B(_1093_),
    .C(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__a21o_1 _4939_ (.A1(_1091_),
    .A2(_1093_),
    .B1(_1097_),
    .X(_1099_));
 sky130_fd_sc_hd__a22oi_1 _4940_ (.A1(_0152_),
    .A2(_0559_),
    .B1(_0153_),
    .B2(_0533_),
    .Y(_1100_));
 sky130_fd_sc_hd__and4_1 _4941_ (.A(_0453_),
    .B(_0152_),
    .C(_0559_),
    .D(_2896_),
    .X(_1101_));
 sky130_fd_sc_hd__nor2_1 _4942_ (.A(_1100_),
    .B(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__nand2_1 _4943_ (.A(_2988_),
    .B(_0490_),
    .Y(_1104_));
 sky130_fd_sc_hd__xnor2_1 _4944_ (.A(_1102_),
    .B(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__nand3_2 _4945_ (.A(_1098_),
    .B(_1099_),
    .C(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__and4_1 _4946_ (.A(\A[0][7] ),
    .B(_0555_),
    .C(_0281_),
    .D(_3014_),
    .X(_1107_));
 sky130_fd_sc_hd__a22o_1 _4947_ (.A1(\A[0][7] ),
    .A2(_0282_),
    .B1(_0241_),
    .B2(_0568_),
    .X(_1108_));
 sky130_fd_sc_hd__and2b_1 _4948_ (.A_N(_1107_),
    .B(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__a21boi_1 _4949_ (.A1(_1089_),
    .A2(_1090_),
    .B1_N(_1088_),
    .Y(_1110_));
 sky130_fd_sc_hd__xnor2_1 _4950_ (.A(_1109_),
    .B(_1110_),
    .Y(_1111_));
 sky130_fd_sc_hd__a22o_1 _4951_ (.A1(_0556_),
    .A2(_0152_),
    .B1(_0559_),
    .B2(_0153_),
    .X(_1112_));
 sky130_fd_sc_hd__nand4_1 _4952_ (.A(_0572_),
    .B(_0152_),
    .C(_0559_),
    .D(_0153_),
    .Y(_1113_));
 sky130_fd_sc_hd__and2_1 _4953_ (.A(\B[0][5] ),
    .B(_0453_),
    .X(_1115_));
 sky130_fd_sc_hd__a21oi_1 _4954_ (.A1(_1112_),
    .A2(_1113_),
    .B1(_1115_),
    .Y(_1116_));
 sky130_fd_sc_hd__and3_1 _4955_ (.A(_1112_),
    .B(_1113_),
    .C(_1115_),
    .X(_1117_));
 sky130_fd_sc_hd__nor2_1 _4956_ (.A(_1116_),
    .B(_1117_),
    .Y(_1118_));
 sky130_fd_sc_hd__nand2_1 _4957_ (.A(_1111_),
    .B(_1118_),
    .Y(_1119_));
 sky130_fd_sc_hd__or2_1 _4958_ (.A(_1111_),
    .B(_1118_),
    .X(_1120_));
 sky130_fd_sc_hd__nand2_1 _4959_ (.A(_1119_),
    .B(_1120_),
    .Y(_1121_));
 sky130_fd_sc_hd__a21oi_1 _4960_ (.A1(_1098_),
    .A2(_1106_),
    .B1(_1121_),
    .Y(_1122_));
 sky130_fd_sc_hd__nand2_1 _4961_ (.A(_1098_),
    .B(_1106_),
    .Y(_1123_));
 sky130_fd_sc_hd__xor2_2 _4962_ (.A(_1121_),
    .B(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__a32o_1 _4963_ (.A1(_0446_),
    .A2(_0085_),
    .A3(_1031_),
    .B1(_1030_),
    .B2(_0964_),
    .X(_1126_));
 sky130_fd_sc_hd__o21ba_1 _4964_ (.A1(_1100_),
    .A2(_1104_),
    .B1_N(_1101_),
    .X(_1127_));
 sky130_fd_sc_hd__and4_1 _4965_ (.A(_2887_),
    .B(\B[0][7] ),
    .C(_0447_),
    .D(_0455_),
    .X(_1128_));
 sky130_fd_sc_hd__a22oi_1 _4966_ (.A1(_2964_),
    .A2(_0489_),
    .B1(_0490_),
    .B2(_2887_),
    .Y(_1129_));
 sky130_fd_sc_hd__or2_1 _4967_ (.A(_1128_),
    .B(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__or2_1 _4968_ (.A(_1127_),
    .B(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__nand2_1 _4969_ (.A(_1127_),
    .B(_1130_),
    .Y(_1132_));
 sky130_fd_sc_hd__and2_1 _4970_ (.A(_1131_),
    .B(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__nand2_1 _4971_ (.A(_1126_),
    .B(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__or2_1 _4972_ (.A(_1126_),
    .B(_1133_),
    .X(_1135_));
 sky130_fd_sc_hd__and2_1 _4973_ (.A(_1134_),
    .B(_1135_),
    .X(_1137_));
 sky130_fd_sc_hd__and2b_1 _4974_ (.A_N(_1124_),
    .B(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__a22o_1 _4975_ (.A1(_0555_),
    .A2(_0152_),
    .B1(_0153_),
    .B2(_0572_),
    .X(_1139_));
 sky130_fd_sc_hd__and4_1 _4976_ (.A(_0555_),
    .B(_0556_),
    .C(_0152_),
    .D(_0153_),
    .X(_1140_));
 sky130_fd_sc_hd__inv_2 _4977_ (.A(_1140_),
    .Y(_1141_));
 sky130_fd_sc_hd__a22oi_1 _4978_ (.A1(_0400_),
    .A2(_0581_),
    .B1(_1139_),
    .B2(_1141_),
    .Y(_1142_));
 sky130_fd_sc_hd__and4b_1 _4979_ (.A_N(_1140_),
    .B(_0581_),
    .C(_2988_),
    .D(_1139_),
    .X(_1143_));
 sky130_fd_sc_hd__nor2_1 _4980_ (.A(_1142_),
    .B(_1143_),
    .Y(_1144_));
 sky130_fd_sc_hd__nand2_1 _4981_ (.A(_0697_),
    .B(_0282_),
    .Y(_1145_));
 sky130_fd_sc_hd__and3_1 _4982_ (.A(_0567_),
    .B(_0241_),
    .C(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__xnor2_1 _4983_ (.A(_1144_),
    .B(_1146_),
    .Y(_1148_));
 sky130_fd_sc_hd__inv_2 _4984_ (.A(_1108_),
    .Y(_1149_));
 sky130_fd_sc_hd__o31ai_1 _4985_ (.A1(_1107_),
    .A2(_1149_),
    .A3(_1110_),
    .B1(_1119_),
    .Y(_1150_));
 sky130_fd_sc_hd__xor2_1 _4986_ (.A(_1148_),
    .B(_1150_),
    .X(_1151_));
 sky130_fd_sc_hd__and4_1 _4987_ (.A(_0572_),
    .B(_0185_),
    .C(_0581_),
    .D(_0186_),
    .X(_1152_));
 sky130_fd_sc_hd__and4_1 _4988_ (.A(_2887_),
    .B(\B[0][7] ),
    .C(_0454_),
    .D(_0453_),
    .X(_1153_));
 sky130_fd_sc_hd__a22oi_1 _4989_ (.A1(_2964_),
    .A2(_0455_),
    .B1(_0533_),
    .B2(_2887_),
    .Y(_1154_));
 sky130_fd_sc_hd__or2_1 _4990_ (.A(_1153_),
    .B(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__o21bai_2 _4991_ (.A1(_1152_),
    .A2(_1117_),
    .B1_N(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__or3b_1 _4992_ (.A(_1152_),
    .B(_1117_),
    .C_N(_1155_),
    .X(_1157_));
 sky130_fd_sc_hd__and2_1 _4993_ (.A(_1156_),
    .B(_1157_),
    .X(_1159_));
 sky130_fd_sc_hd__or2_1 _4994_ (.A(_1159_),
    .B(_1128_),
    .X(_1160_));
 sky130_fd_sc_hd__nand2_1 _4995_ (.A(_1159_),
    .B(_1128_),
    .Y(_1161_));
 sky130_fd_sc_hd__nand2_1 _4996_ (.A(_1160_),
    .B(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__xor2_1 _4997_ (.A(_1151_),
    .B(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__o21a_1 _4998_ (.A1(_1122_),
    .A2(_1138_),
    .B1(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__nor3_1 _4999_ (.A(_1163_),
    .B(_1122_),
    .C(_1138_),
    .Y(_1165_));
 sky130_fd_sc_hd__nor2_1 _5000_ (.A(_1164_),
    .B(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__nand2_1 _5001_ (.A(_1055_),
    .B(_1058_),
    .Y(_1167_));
 sky130_fd_sc_hd__o21a_1 _5002_ (.A1(_1050_),
    .A2(_1060_),
    .B1(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__a22oi_1 _5003_ (.A1(_0159_),
    .A2(_0500_),
    .B1(_0160_),
    .B2(_0502_),
    .Y(_1170_));
 sky130_fd_sc_hd__and4_1 _5004_ (.A(_0159_),
    .B(_0502_),
    .C(_0430_),
    .D(_2917_),
    .X(_1171_));
 sky130_fd_sc_hd__nor2_1 _5005_ (.A(_1170_),
    .B(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__nand2_1 _5006_ (.A(_2921_),
    .B(_0506_),
    .Y(_1173_));
 sky130_fd_sc_hd__xnor2_1 _5007_ (.A(_1172_),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__a22oi_1 _5008_ (.A1(\A[1][7] ),
    .A2(_0220_),
    .B1(_3001_),
    .B2(_0443_),
    .Y(_1175_));
 sky130_fd_sc_hd__and4_1 _5009_ (.A(\A[1][7] ),
    .B(_0422_),
    .C(_0220_),
    .D(\B[2][3] ),
    .X(_1176_));
 sky130_fd_sc_hd__or2_1 _5010_ (.A(_1175_),
    .B(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__and4_1 _5011_ (.A(\A[1][7] ),
    .B(_0443_),
    .C(_0221_),
    .D(_0220_),
    .X(_1178_));
 sky130_fd_sc_hd__a31o_1 _5012_ (.A1(_0502_),
    .A2(_3001_),
    .A3(_1052_),
    .B1(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__xnor2_1 _5013_ (.A(_1177_),
    .B(_1179_),
    .Y(_1181_));
 sky130_fd_sc_hd__nand2_1 _5014_ (.A(_1174_),
    .B(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__or2_1 _5015_ (.A(_1174_),
    .B(_1181_),
    .X(_1183_));
 sky130_fd_sc_hd__nand2_1 _5016_ (.A(_1182_),
    .B(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__a21oi_1 _5017_ (.A1(_1131_),
    .A2(_1134_),
    .B1(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__and3_1 _5018_ (.A(_1131_),
    .B(_1134_),
    .C(_1184_),
    .X(_1186_));
 sky130_fd_sc_hd__nor2_1 _5019_ (.A(_1185_),
    .B(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__xnor2_1 _5020_ (.A(_1168_),
    .B(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__xnor2_1 _5021_ (.A(_1166_),
    .B(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__xnor2_1 _5022_ (.A(_1078_),
    .B(_1080_),
    .Y(_1190_));
 sky130_fd_sc_hd__xnor2_2 _5023_ (.A(_1124_),
    .B(_1137_),
    .Y(_1192_));
 sky130_fd_sc_hd__xor2_2 _5024_ (.A(_1041_),
    .B(_1042_),
    .X(_1193_));
 sky130_fd_sc_hd__a21o_1 _5025_ (.A1(_1098_),
    .A2(_1099_),
    .B1(_1105_),
    .X(_1194_));
 sky130_fd_sc_hd__o2bb2a_1 _5026_ (.A1_N(_0400_),
    .A2_N(_0531_),
    .B1(_1035_),
    .B2(_1036_),
    .X(_1195_));
 sky130_fd_sc_hd__nor2_1 _5027_ (.A(_1038_),
    .B(_1195_),
    .Y(_1196_));
 sky130_fd_sc_hd__or3_1 _5028_ (.A(_1096_),
    .B(_1094_),
    .C(_1095_),
    .X(_1197_));
 sky130_fd_sc_hd__o21ai_1 _5029_ (.A1(_1096_),
    .A2(_1094_),
    .B1(_1095_),
    .Y(_1198_));
 sky130_fd_sc_hd__nand2_1 _5030_ (.A(_0241_),
    .B(_0453_),
    .Y(_1199_));
 sky130_fd_sc_hd__a22oi_2 _5031_ (.A1(_0556_),
    .A2(_0279_),
    .B1(_0281_),
    .B2(_0559_),
    .Y(_1200_));
 sky130_fd_sc_hd__and4_1 _5032_ (.A(_0556_),
    .B(_3046_),
    .C(_0281_),
    .D(_0493_),
    .X(_1201_));
 sky130_fd_sc_hd__o21bai_1 _5033_ (.A1(_1199_),
    .A2(_1200_),
    .B1_N(_1201_),
    .Y(_1203_));
 sky130_fd_sc_hd__a21o_1 _5034_ (.A1(_1197_),
    .A2(_1198_),
    .B1(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__nand3_1 _5035_ (.A(_1197_),
    .B(_1198_),
    .C(_1203_),
    .Y(_1205_));
 sky130_fd_sc_hd__a21bo_1 _5036_ (.A1(_1196_),
    .A2(_1204_),
    .B1_N(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__a21o_1 _5037_ (.A1(_1106_),
    .A2(_1194_),
    .B1(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__nand3_2 _5038_ (.A(_1106_),
    .B(_1194_),
    .C(_1206_),
    .Y(_1208_));
 sky130_fd_sc_hd__a21boi_2 _5039_ (.A1(_1193_),
    .A2(_1207_),
    .B1_N(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__xnor2_1 _5040_ (.A(_1192_),
    .B(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__or2b_1 _5041_ (.A(_1209_),
    .B_N(_1192_),
    .X(_1211_));
 sky130_fd_sc_hd__a21bo_1 _5042_ (.A1(_1190_),
    .A2(_1210_),
    .B1_N(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__and2b_1 _5043_ (.A_N(_1189_),
    .B(_1212_),
    .X(_1214_));
 sky130_fd_sc_hd__nand2_1 _5044_ (.A(_2886_),
    .B(_0421_),
    .Y(_1215_));
 sky130_fd_sc_hd__xor2_1 _5045_ (.A(_1086_),
    .B(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__xor2_1 _5046_ (.A(_1189_),
    .B(_1212_),
    .X(_1217_));
 sky130_fd_sc_hd__nor2_1 _5047_ (.A(_1216_),
    .B(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__nand2_1 _5048_ (.A(_0567_),
    .B(_0185_),
    .Y(_1219_));
 sky130_fd_sc_hd__nand2_1 _5049_ (.A(_0568_),
    .B(_0186_),
    .Y(_1220_));
 sky130_fd_sc_hd__and4_1 _5050_ (.A(_0567_),
    .B(_0568_),
    .C(_0185_),
    .D(_0186_),
    .X(_1221_));
 sky130_fd_sc_hd__a21oi_1 _5051_ (.A1(_1219_),
    .A2(_1220_),
    .B1(_1221_),
    .Y(_1222_));
 sky130_fd_sc_hd__nand2_1 _5052_ (.A(_0400_),
    .B(_0573_),
    .Y(_1223_));
 sky130_fd_sc_hd__xnor2_1 _5053_ (.A(_1222_),
    .B(_1223_),
    .Y(_1225_));
 sky130_fd_sc_hd__a21oi_1 _5054_ (.A1(_1144_),
    .A2(_1146_),
    .B1(_1107_),
    .Y(_1226_));
 sky130_fd_sc_hd__xnor2_1 _5055_ (.A(_1225_),
    .B(_1226_),
    .Y(_1227_));
 sky130_fd_sc_hd__or2_1 _5056_ (.A(_1140_),
    .B(_1143_),
    .X(_1228_));
 sky130_fd_sc_hd__clkbuf_4 _5057_ (.A(_2964_),
    .X(_1229_));
 sky130_fd_sc_hd__a22o_1 _5058_ (.A1(_1229_),
    .A2(_0533_),
    .B1(_0581_),
    .B2(_2888_),
    .X(_1230_));
 sky130_fd_sc_hd__and3_1 _5059_ (.A(_2888_),
    .B(_2964_),
    .C(_0581_),
    .X(_1231_));
 sky130_fd_sc_hd__nand2_1 _5060_ (.A(_0533_),
    .B(_1231_),
    .Y(_1232_));
 sky130_fd_sc_hd__nand2_1 _5061_ (.A(_1230_),
    .B(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__xor2_2 _5062_ (.A(_1228_),
    .B(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__xor2_2 _5063_ (.A(_1234_),
    .B(_1153_),
    .X(_1236_));
 sky130_fd_sc_hd__xnor2_2 _5064_ (.A(_1227_),
    .B(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__or2b_1 _5065_ (.A(_1148_),
    .B_N(_1150_),
    .X(_1238_));
 sky130_fd_sc_hd__o21ai_2 _5066_ (.A1(_1151_),
    .A2(_1162_),
    .B1(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__xor2_1 _5067_ (.A(_1237_),
    .B(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__or2b_1 _5068_ (.A(_1177_),
    .B_N(_1179_),
    .X(_1241_));
 sky130_fd_sc_hd__nand2_1 _5069_ (.A(_1241_),
    .B(_1182_),
    .Y(_1242_));
 sky130_fd_sc_hd__a22oi_1 _5070_ (.A1(_0159_),
    .A2(_0502_),
    .B1(_0160_),
    .B2(_0443_),
    .Y(_1243_));
 sky130_fd_sc_hd__and2_1 _5071_ (.A(_2916_),
    .B(_0422_),
    .X(_1244_));
 sky130_fd_sc_hd__and3_1 _5072_ (.A(_0502_),
    .B(_0160_),
    .C(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__nor2_1 _5073_ (.A(_1243_),
    .B(_1245_),
    .Y(_1247_));
 sky130_fd_sc_hd__nand2_1 _5074_ (.A(_2921_),
    .B(_0500_),
    .Y(_1248_));
 sky130_fd_sc_hd__xnor2_1 _5075_ (.A(_1247_),
    .B(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__nand2_1 _5076_ (.A(_0546_),
    .B(_0294_),
    .Y(_1250_));
 sky130_fd_sc_hd__and3_1 _5077_ (.A(_0446_),
    .B(_3002_),
    .C(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__xnor2_1 _5078_ (.A(_1249_),
    .B(_1251_),
    .Y(_1252_));
 sky130_fd_sc_hd__a21oi_1 _5079_ (.A1(_1156_),
    .A2(_1161_),
    .B1(_1252_),
    .Y(_1253_));
 sky130_fd_sc_hd__and3_1 _5080_ (.A(_1156_),
    .B(_1161_),
    .C(_1252_),
    .X(_1254_));
 sky130_fd_sc_hd__or2_1 _5081_ (.A(_1253_),
    .B(_1254_),
    .X(_1255_));
 sky130_fd_sc_hd__xnor2_1 _5082_ (.A(_1242_),
    .B(_1255_),
    .Y(_1256_));
 sky130_fd_sc_hd__nand2_1 _5083_ (.A(_1240_),
    .B(_1256_),
    .Y(_1258_));
 sky130_fd_sc_hd__or2_1 _5084_ (.A(_1240_),
    .B(_1256_),
    .X(_1259_));
 sky130_fd_sc_hd__nand2_1 _5085_ (.A(_1258_),
    .B(_1259_),
    .Y(_1260_));
 sky130_fd_sc_hd__a21oi_1 _5086_ (.A1(_1166_),
    .A2(_1188_),
    .B1(_1164_),
    .Y(_1261_));
 sky130_fd_sc_hd__xnor2_1 _5087_ (.A(_1260_),
    .B(_1261_),
    .Y(_1262_));
 sky130_fd_sc_hd__and2b_1 _5088_ (.A_N(_1168_),
    .B(_1187_),
    .X(_1263_));
 sky130_fd_sc_hd__o21ba_1 _5089_ (.A1(_1170_),
    .A2(_1173_),
    .B1_N(_1171_),
    .X(_1264_));
 sky130_fd_sc_hd__o21ba_1 _5090_ (.A1(_1185_),
    .A2(_1263_),
    .B1_N(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__or3b_1 _5091_ (.A(_1185_),
    .B(_1263_),
    .C_N(_1264_),
    .X(_1266_));
 sky130_fd_sc_hd__and2b_1 _5092_ (.A_N(_1265_),
    .B(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__nand2_1 _5093_ (.A(_2886_),
    .B(_0506_),
    .Y(_1269_));
 sky130_fd_sc_hd__xor2_1 _5094_ (.A(_1267_),
    .B(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__xor2_1 _5095_ (.A(_1262_),
    .B(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__o21ai_1 _5096_ (.A1(_1214_),
    .A2(_1218_),
    .B1(_1271_),
    .Y(_1272_));
 sky130_fd_sc_hd__or3_1 _5097_ (.A(_1271_),
    .B(_1214_),
    .C(_1218_),
    .X(_1273_));
 sky130_fd_sc_hd__and2_1 _5098_ (.A(_1272_),
    .B(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__xnor2_2 _5099_ (.A(_1087_),
    .B(_1274_),
    .Y(_1275_));
 sky130_fd_sc_hd__a22oi_1 _5100_ (.A1(_0490_),
    .A2(_0185_),
    .B1(_0186_),
    .B2(_0489_),
    .Y(_1276_));
 sky130_fd_sc_hd__and4_1 _5101_ (.A(_0489_),
    .B(_0455_),
    .C(_0152_),
    .D(_0153_),
    .X(_1277_));
 sky130_fd_sc_hd__nor2_1 _5102_ (.A(_1276_),
    .B(_1277_),
    .Y(_1278_));
 sky130_fd_sc_hd__a31o_1 _5103_ (.A1(_0400_),
    .A2(_0964_),
    .A3(_1278_),
    .B1(_1277_),
    .X(_1280_));
 sky130_fd_sc_hd__a22oi_1 _5104_ (.A1(_2888_),
    .A2(_0726_),
    .B1(_0085_),
    .B2(_0546_),
    .Y(_1281_));
 sky130_fd_sc_hd__nor2_1 _5105_ (.A(_1042_),
    .B(_1281_),
    .Y(_1282_));
 sky130_fd_sc_hd__nand2_2 _5106_ (.A(_1280_),
    .B(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__xnor2_1 _5107_ (.A(_1067_),
    .B(_1076_),
    .Y(_1284_));
 sky130_fd_sc_hd__nor2_1 _5108_ (.A(_1283_),
    .B(_1284_),
    .Y(_1285_));
 sky130_fd_sc_hd__a22oi_1 _5109_ (.A1(_0159_),
    .A2(_0719_),
    .B1(_0420_),
    .B2(_0160_),
    .Y(_1286_));
 sky130_fd_sc_hd__and4_1 _5110_ (.A(_0159_),
    .B(_0476_),
    .C(_0420_),
    .D(_0160_),
    .X(_1287_));
 sky130_fd_sc_hd__nor2_1 _5111_ (.A(_1286_),
    .B(_1287_),
    .Y(_1288_));
 sky130_fd_sc_hd__nand2_1 _5112_ (.A(_2921_),
    .B(_0810_),
    .Y(_1289_));
 sky130_fd_sc_hd__xnor2_1 _5113_ (.A(_1288_),
    .B(_1289_),
    .Y(_1291_));
 sky130_fd_sc_hd__o2bb2a_1 _5114_ (.A1_N(_0472_),
    .A2_N(_3001_),
    .B1(_1072_),
    .B2(_1073_),
    .X(_1292_));
 sky130_fd_sc_hd__nor2_1 _5115_ (.A(_1074_),
    .B(_1292_),
    .Y(_1293_));
 sky130_fd_sc_hd__and4_1 _5116_ (.A(_0221_),
    .B(_0220_),
    .C(_0436_),
    .D(_0430_),
    .X(_1294_));
 sky130_fd_sc_hd__a22oi_1 _5117_ (.A1(_0294_),
    .A2(_0472_),
    .B1(_0500_),
    .B2(_0293_),
    .Y(_1295_));
 sky130_fd_sc_hd__and4bb_1 _5118_ (.A_N(_1294_),
    .B_N(_1295_),
    .C(_0420_),
    .D(_3001_),
    .X(_1296_));
 sky130_fd_sc_hd__nor2_1 _5119_ (.A(_1294_),
    .B(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__xnor2_1 _5120_ (.A(_1293_),
    .B(_1297_),
    .Y(_1298_));
 sky130_fd_sc_hd__and2b_1 _5121_ (.A_N(_1297_),
    .B(_1293_),
    .X(_1299_));
 sky130_fd_sc_hd__a21o_1 _5122_ (.A1(_1291_),
    .A2(_1298_),
    .B1(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__xor2_1 _5123_ (.A(_1283_),
    .B(_1284_),
    .X(_1302_));
 sky130_fd_sc_hd__and2_1 _5124_ (.A(_1300_),
    .B(_1302_),
    .X(_1303_));
 sky130_fd_sc_hd__o21ba_1 _5125_ (.A1(_1063_),
    .A2(_1066_),
    .B1_N(_1064_),
    .X(_1304_));
 sky130_fd_sc_hd__o21ba_1 _5126_ (.A1(_1285_),
    .A2(_1303_),
    .B1_N(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__or3b_1 _5127_ (.A(_1285_),
    .B(_1303_),
    .C_N(_1304_),
    .X(_1306_));
 sky130_fd_sc_hd__and2b_1 _5128_ (.A_N(_1305_),
    .B(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__a31o_1 _5129_ (.A1(_1029_),
    .A2(_0720_),
    .A3(_1307_),
    .B1(_1305_),
    .X(_1308_));
 sky130_fd_sc_hd__xor2_1 _5130_ (.A(_1216_),
    .B(_1217_),
    .X(_1309_));
 sky130_fd_sc_hd__nand2_1 _5131_ (.A(_2886_),
    .B(_0720_),
    .Y(_1310_));
 sky130_fd_sc_hd__xor2_1 _5132_ (.A(_1307_),
    .B(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__xnor2_1 _5133_ (.A(_1190_),
    .B(_1210_),
    .Y(_1313_));
 sky130_fd_sc_hd__nand3_1 _5134_ (.A(_1205_),
    .B(_1196_),
    .C(_1204_),
    .Y(_1314_));
 sky130_fd_sc_hd__a21o_1 _5135_ (.A1(_1205_),
    .A2(_1204_),
    .B1(_1196_),
    .X(_1315_));
 sky130_fd_sc_hd__nand2_1 _5136_ (.A(_2988_),
    .B(_0726_),
    .Y(_1316_));
 sky130_fd_sc_hd__xnor2_1 _5137_ (.A(_1278_),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__or3_1 _5138_ (.A(_1201_),
    .B(_1199_),
    .C(_1200_),
    .X(_1318_));
 sky130_fd_sc_hd__o21ai_1 _5139_ (.A1(_1201_),
    .A2(_1200_),
    .B1(_1199_),
    .Y(_1319_));
 sky130_fd_sc_hd__nand2_1 _5140_ (.A(_0455_),
    .B(_3014_),
    .Y(_1320_));
 sky130_fd_sc_hd__a22oi_2 _5141_ (.A1(_0281_),
    .A2(_0453_),
    .B1(_0559_),
    .B2(_0279_),
    .Y(_1321_));
 sky130_fd_sc_hd__and4_1 _5142_ (.A(_0279_),
    .B(_0281_),
    .C(_0457_),
    .D(_0493_),
    .X(_1322_));
 sky130_fd_sc_hd__o21bai_1 _5143_ (.A1(_1320_),
    .A2(_1321_),
    .B1_N(_1322_),
    .Y(_1324_));
 sky130_fd_sc_hd__a21o_1 _5144_ (.A1(_1318_),
    .A2(_1319_),
    .B1(_1324_),
    .X(_1325_));
 sky130_fd_sc_hd__nand3_1 _5145_ (.A(_1318_),
    .B(_1319_),
    .C(_1324_),
    .Y(_1326_));
 sky130_fd_sc_hd__a21bo_1 _5146_ (.A1(_1317_),
    .A2(_1325_),
    .B1_N(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__nand3_4 _5147_ (.A(_1314_),
    .B(_1315_),
    .C(_1327_),
    .Y(_1328_));
 sky130_fd_sc_hd__or2_1 _5148_ (.A(_1280_),
    .B(_1282_),
    .X(_1329_));
 sky130_fd_sc_hd__and2_1 _5149_ (.A(_1283_),
    .B(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__a21o_1 _5150_ (.A1(_1314_),
    .A2(_1315_),
    .B1(_1327_),
    .X(_1331_));
 sky130_fd_sc_hd__nand3_4 _5151_ (.A(_1328_),
    .B(_1330_),
    .C(_1331_),
    .Y(_1332_));
 sky130_fd_sc_hd__and3_1 _5152_ (.A(_1208_),
    .B(_1193_),
    .C(_1207_),
    .X(_1333_));
 sky130_fd_sc_hd__a21oi_2 _5153_ (.A1(_1208_),
    .A2(_1207_),
    .B1(_1193_),
    .Y(_1335_));
 sky130_fd_sc_hd__a211o_1 _5154_ (.A1(_1328_),
    .A2(_1332_),
    .B1(_1333_),
    .C1(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__xnor2_1 _5155_ (.A(_1300_),
    .B(_1302_),
    .Y(_1337_));
 sky130_fd_sc_hd__o211ai_4 _5156_ (.A1(_1333_),
    .A2(_1335_),
    .B1(_1328_),
    .C1(_1332_),
    .Y(_1338_));
 sky130_fd_sc_hd__nand3b_1 _5157_ (.A_N(_1337_),
    .B(_1338_),
    .C(_1336_),
    .Y(_1339_));
 sky130_fd_sc_hd__nand2_1 _5158_ (.A(_1336_),
    .B(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__xor2_1 _5159_ (.A(_1313_),
    .B(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__or2b_1 _5160_ (.A(_1313_),
    .B_N(_1340_),
    .X(_1342_));
 sky130_fd_sc_hd__o21a_1 _5161_ (.A1(_1311_),
    .A2(_1341_),
    .B1(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__xnor2_1 _5162_ (.A(_1309_),
    .B(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__or2b_1 _5163_ (.A(_1343_),
    .B_N(_1309_),
    .X(_1346_));
 sky130_fd_sc_hd__a21boi_1 _5164_ (.A1(_1308_),
    .A2(_1344_),
    .B1_N(_1346_),
    .Y(_1347_));
 sky130_fd_sc_hd__or2_2 _5165_ (.A(_1275_),
    .B(_1347_),
    .X(_1348_));
 sky130_fd_sc_hd__xnor2_2 _5166_ (.A(_1275_),
    .B(_1347_),
    .Y(_1349_));
 sky130_fd_sc_hd__xnor2_1 _5167_ (.A(_1308_),
    .B(_1344_),
    .Y(_1350_));
 sky130_fd_sc_hd__nand3_1 _5168_ (.A(_1326_),
    .B(_1317_),
    .C(_1325_),
    .Y(_1351_));
 sky130_fd_sc_hd__a21o_1 _5169_ (.A1(_1326_),
    .A2(_1325_),
    .B1(_1317_),
    .X(_1352_));
 sky130_fd_sc_hd__and4_1 _5170_ (.A(_0444_),
    .B(_0489_),
    .C(_0185_),
    .D(_0186_),
    .X(_1353_));
 sky130_fd_sc_hd__a22oi_1 _5171_ (.A1(_0531_),
    .A2(_0185_),
    .B1(_0186_),
    .B2(_0726_),
    .Y(_1354_));
 sky130_fd_sc_hd__nor2_1 _5172_ (.A(_1353_),
    .B(_1354_),
    .Y(_1355_));
 sky130_fd_sc_hd__or3_1 _5173_ (.A(_1322_),
    .B(_1320_),
    .C(_1321_),
    .X(_1357_));
 sky130_fd_sc_hd__o21ai_1 _5174_ (.A1(_1322_),
    .A2(_1321_),
    .B1(_1320_),
    .Y(_1358_));
 sky130_fd_sc_hd__nand2_1 _5175_ (.A(_0447_),
    .B(_3014_),
    .Y(_1359_));
 sky130_fd_sc_hd__a22oi_2 _5176_ (.A1(_0281_),
    .A2(_0454_),
    .B1(_0457_),
    .B2(_0279_),
    .Y(_1360_));
 sky130_fd_sc_hd__and4_1 _5177_ (.A(_3046_),
    .B(_3015_),
    .C(_0454_),
    .D(_0457_),
    .X(_1361_));
 sky130_fd_sc_hd__o21bai_1 _5178_ (.A1(_1359_),
    .A2(_1360_),
    .B1_N(_1361_),
    .Y(_1362_));
 sky130_fd_sc_hd__a21o_1 _5179_ (.A1(_1357_),
    .A2(_1358_),
    .B1(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__nand3_1 _5180_ (.A(_1357_),
    .B(_1358_),
    .C(_1362_),
    .Y(_1364_));
 sky130_fd_sc_hd__a21bo_1 _5181_ (.A1(_1355_),
    .A2(_1363_),
    .B1_N(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__and3_2 _5182_ (.A(_1351_),
    .B(_1352_),
    .C(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__nand3_2 _5183_ (.A(_0684_),
    .B(_0085_),
    .C(_1353_),
    .Y(_1368_));
 sky130_fd_sc_hd__a21o_1 _5184_ (.A1(_0684_),
    .A2(_0085_),
    .B1(_1353_),
    .X(_1369_));
 sky130_fd_sc_hd__nand2_1 _5185_ (.A(_1368_),
    .B(_1369_),
    .Y(_1370_));
 sky130_fd_sc_hd__a21oi_2 _5186_ (.A1(_1351_),
    .A2(_1352_),
    .B1(_1365_),
    .Y(_1371_));
 sky130_fd_sc_hd__nor3_4 _5187_ (.A(_1366_),
    .B(_1370_),
    .C(_1371_),
    .Y(_1372_));
 sky130_fd_sc_hd__a21o_1 _5188_ (.A1(_1328_),
    .A2(_1331_),
    .B1(_1330_),
    .X(_1373_));
 sky130_fd_sc_hd__o211a_2 _5189_ (.A1(_1366_),
    .A2(_1372_),
    .B1(_1332_),
    .C1(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__o2bb2a_1 _5190_ (.A1_N(_0421_),
    .A2_N(_3002_),
    .B1(_1294_),
    .B2(_1295_),
    .X(_1375_));
 sky130_fd_sc_hd__and4_1 _5191_ (.A(_0221_),
    .B(_0419_),
    .C(_0220_),
    .D(_0436_),
    .X(_1376_));
 sky130_fd_sc_hd__a22oi_1 _5192_ (.A1(_0420_),
    .A2(_0294_),
    .B1(_0472_),
    .B2(_0293_),
    .Y(_1377_));
 sky130_fd_sc_hd__and4bb_1 _5193_ (.A_N(_1376_),
    .B_N(_1377_),
    .C(_0719_),
    .D(_3001_),
    .X(_1379_));
 sky130_fd_sc_hd__nor2_1 _5194_ (.A(_1376_),
    .B(_1379_),
    .Y(_1380_));
 sky130_fd_sc_hd__or3_1 _5195_ (.A(_1296_),
    .B(_1375_),
    .C(_1380_),
    .X(_1381_));
 sky130_fd_sc_hd__nor2_1 _5196_ (.A(_1296_),
    .B(_1375_),
    .Y(_1382_));
 sky130_fd_sc_hd__xnor2_1 _5197_ (.A(_1382_),
    .B(_1380_),
    .Y(_1383_));
 sky130_fd_sc_hd__a22oi_1 _5198_ (.A1(_0378_),
    .A2(\A[1][0] ),
    .B1(_0719_),
    .B2(_0229_),
    .Y(_1384_));
 sky130_fd_sc_hd__and4_1 _5199_ (.A(_0378_),
    .B(\A[1][0] ),
    .C(_0719_),
    .D(_0160_),
    .X(_1385_));
 sky130_fd_sc_hd__or2_1 _5200_ (.A(_1384_),
    .B(_1385_),
    .X(_1386_));
 sky130_fd_sc_hd__inv_2 _5201_ (.A(_1386_),
    .Y(_1387_));
 sky130_fd_sc_hd__nand2_1 _5202_ (.A(_1383_),
    .B(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__xnor2_1 _5203_ (.A(_1291_),
    .B(_1298_),
    .Y(_1390_));
 sky130_fd_sc_hd__xnor2_1 _5204_ (.A(_1368_),
    .B(_1390_),
    .Y(_1391_));
 sky130_fd_sc_hd__a21oi_2 _5205_ (.A1(_1381_),
    .A2(_1388_),
    .B1(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__and3_1 _5206_ (.A(_1381_),
    .B(_1388_),
    .C(_1391_),
    .X(_1393_));
 sky130_fd_sc_hd__a211oi_4 _5207_ (.A1(_1332_),
    .A2(_1373_),
    .B1(_1366_),
    .C1(_1372_),
    .Y(_1394_));
 sky130_fd_sc_hd__nor4_1 _5208_ (.A(_1374_),
    .B(_1392_),
    .C(_1393_),
    .D(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__a21bo_1 _5209_ (.A1(_1336_),
    .A2(_1338_),
    .B1_N(_1337_),
    .X(_1396_));
 sky130_fd_sc_hd__o211ai_2 _5210_ (.A1(_1374_),
    .A2(_1395_),
    .B1(_1339_),
    .C1(_1396_),
    .Y(_1397_));
 sky130_fd_sc_hd__nor2_1 _5211_ (.A(_1368_),
    .B(_1390_),
    .Y(_1398_));
 sky130_fd_sc_hd__o21ba_1 _5212_ (.A1(_1286_),
    .A2(_1289_),
    .B1_N(_1287_),
    .X(_1399_));
 sky130_fd_sc_hd__o21ba_1 _5213_ (.A1(_1398_),
    .A2(_1392_),
    .B1_N(_1399_),
    .X(_1401_));
 sky130_fd_sc_hd__or3b_1 _5214_ (.A(_1398_),
    .B(_1392_),
    .C_N(_1399_),
    .X(_1402_));
 sky130_fd_sc_hd__and2b_1 _5215_ (.A_N(_1401_),
    .B(_1402_),
    .X(_1403_));
 sky130_fd_sc_hd__nand2_1 _5216_ (.A(_2886_),
    .B(_0899_),
    .Y(_1404_));
 sky130_fd_sc_hd__xor2_1 _5217_ (.A(_1403_),
    .B(_1404_),
    .X(_1405_));
 sky130_fd_sc_hd__a211o_1 _5218_ (.A1(_1339_),
    .A2(_1396_),
    .B1(_1374_),
    .C1(_1395_),
    .X(_1406_));
 sky130_fd_sc_hd__nand2_1 _5219_ (.A(_1397_),
    .B(_1406_),
    .Y(_1407_));
 sky130_fd_sc_hd__or2_1 _5220_ (.A(_1405_),
    .B(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__xnor2_1 _5221_ (.A(_1311_),
    .B(_1341_),
    .Y(_1409_));
 sky130_fd_sc_hd__a21o_1 _5222_ (.A1(_1397_),
    .A2(_1408_),
    .B1(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__a21oi_1 _5223_ (.A1(_1397_),
    .A2(_1408_),
    .B1(_1409_),
    .Y(_1412_));
 sky130_fd_sc_hd__a31oi_2 _5224_ (.A1(_1029_),
    .A2(_0899_),
    .A3(_1403_),
    .B1(_1401_),
    .Y(_1413_));
 sky130_fd_sc_hd__and3_1 _5225_ (.A(_1409_),
    .B(_1397_),
    .C(_1408_),
    .X(_1414_));
 sky130_fd_sc_hd__or3_1 _5226_ (.A(_1412_),
    .B(_1413_),
    .C(_1414_),
    .X(_1415_));
 sky130_fd_sc_hd__and3_1 _5227_ (.A(_1350_),
    .B(_1410_),
    .C(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__nor2_1 _5228_ (.A(_1412_),
    .B(_1414_),
    .Y(_1417_));
 sky130_fd_sc_hd__xnor2_1 _5229_ (.A(_1413_),
    .B(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__o2bb2a_1 _5230_ (.A1_N(_0719_),
    .A2_N(_3002_),
    .B1(_1376_),
    .B2(_1377_),
    .X(_1419_));
 sky130_fd_sc_hd__and4_1 _5231_ (.A(_0476_),
    .B(_0221_),
    .C(_0419_),
    .D(_0220_),
    .X(_1420_));
 sky130_fd_sc_hd__a22oi_1 _5232_ (.A1(_0293_),
    .A2(_0420_),
    .B1(_0294_),
    .B2(_0476_),
    .Y(_1421_));
 sky130_fd_sc_hd__and4bb_1 _5233_ (.A_N(_1420_),
    .B_N(_1421_),
    .C(\A[1][0] ),
    .D(_3001_),
    .X(_1423_));
 sky130_fd_sc_hd__nor2_1 _5234_ (.A(_1420_),
    .B(_1423_),
    .Y(_1424_));
 sky130_fd_sc_hd__or3_1 _5235_ (.A(_1379_),
    .B(_1419_),
    .C(_1424_),
    .X(_1425_));
 sky130_fd_sc_hd__nand2_1 _5236_ (.A(_0810_),
    .B(_0229_),
    .Y(_1426_));
 sky130_fd_sc_hd__nor2_1 _5237_ (.A(_1379_),
    .B(_1419_),
    .Y(_1427_));
 sky130_fd_sc_hd__xnor2_1 _5238_ (.A(_1427_),
    .B(_1424_),
    .Y(_1428_));
 sky130_fd_sc_hd__or2b_1 _5239_ (.A(_1426_),
    .B_N(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__xnor2_1 _5240_ (.A(_1383_),
    .B(_1387_),
    .Y(_1430_));
 sky130_fd_sc_hd__a21oi_1 _5241_ (.A1(_1425_),
    .A2(_1429_),
    .B1(_1430_),
    .Y(_1431_));
 sky130_fd_sc_hd__and2_1 _5242_ (.A(_1385_),
    .B(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__xor2_1 _5243_ (.A(_1405_),
    .B(_1407_),
    .X(_1434_));
 sky130_fd_sc_hd__nand3_1 _5244_ (.A(_1364_),
    .B(_1355_),
    .C(_1363_),
    .Y(_1435_));
 sky130_fd_sc_hd__a21o_1 _5245_ (.A1(_1364_),
    .A2(_1363_),
    .B1(_1355_),
    .X(_1436_));
 sky130_fd_sc_hd__nand2_1 _5246_ (.A(_0964_),
    .B(_0185_),
    .Y(_1437_));
 sky130_fd_sc_hd__or3_1 _5247_ (.A(_1361_),
    .B(_1359_),
    .C(_1360_),
    .X(_1438_));
 sky130_fd_sc_hd__o21ai_1 _5248_ (.A1(_1361_),
    .A2(_1360_),
    .B1(_1359_),
    .Y(_1439_));
 sky130_fd_sc_hd__a22o_1 _5249_ (.A1(_0447_),
    .A2(_0281_),
    .B1(_0455_),
    .B2(_0279_),
    .X(_1440_));
 sky130_fd_sc_hd__and4_1 _5250_ (.A(_0279_),
    .B(_0447_),
    .C(_0281_),
    .D(_0454_),
    .X(_1441_));
 sky130_fd_sc_hd__a31o_1 _5251_ (.A1(_0444_),
    .A2(_0241_),
    .A3(_1440_),
    .B1(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__a21oi_2 _5252_ (.A1(_1438_),
    .A2(_1439_),
    .B1(_1442_),
    .Y(_1443_));
 sky130_fd_sc_hd__and3_1 _5253_ (.A(_1438_),
    .B(_1439_),
    .C(_1442_),
    .X(_1445_));
 sky130_fd_sc_hd__o21bai_2 _5254_ (.A1(_1437_),
    .A2(_1443_),
    .B1_N(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__nand3_4 _5255_ (.A(_1435_),
    .B(_1436_),
    .C(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__a21o_1 _5256_ (.A1(_1435_),
    .A2(_1436_),
    .B1(_1446_),
    .X(_1448_));
 sky130_fd_sc_hd__nand4_2 _5257_ (.A(_0342_),
    .B(_0671_),
    .C(_1447_),
    .D(_1448_),
    .Y(_1449_));
 sky130_fd_sc_hd__o21a_1 _5258_ (.A1(_1366_),
    .A2(_1371_),
    .B1(_1370_),
    .X(_1450_));
 sky130_fd_sc_hd__a211oi_2 _5259_ (.A1(_1447_),
    .A2(_1449_),
    .B1(_1372_),
    .C1(_1450_),
    .Y(_1451_));
 sky130_fd_sc_hd__and3_1 _5260_ (.A(_1430_),
    .B(_1425_),
    .C(_1429_),
    .X(_1452_));
 sky130_fd_sc_hd__or2_1 _5261_ (.A(_1431_),
    .B(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__o211a_1 _5262_ (.A1(_1372_),
    .A2(_1450_),
    .B1(_1447_),
    .C1(_1449_),
    .X(_1454_));
 sky130_fd_sc_hd__nor3_2 _5263_ (.A(_1451_),
    .B(_1453_),
    .C(_1454_),
    .Y(_1456_));
 sky130_fd_sc_hd__or4_1 _5264_ (.A(_1374_),
    .B(_1392_),
    .C(_1393_),
    .D(_1394_),
    .X(_1457_));
 sky130_fd_sc_hd__o22ai_1 _5265_ (.A1(_1392_),
    .A2(_1393_),
    .B1(_1394_),
    .B2(_1374_),
    .Y(_1458_));
 sky130_fd_sc_hd__o211a_1 _5266_ (.A1(_1451_),
    .A2(_1456_),
    .B1(_1457_),
    .C1(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__nor2_1 _5267_ (.A(_1385_),
    .B(_1431_),
    .Y(_1460_));
 sky130_fd_sc_hd__or2_1 _5268_ (.A(_1432_),
    .B(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__a211oi_1 _5269_ (.A1(_1457_),
    .A2(_1458_),
    .B1(_1451_),
    .C1(_1456_),
    .Y(_1462_));
 sky130_fd_sc_hd__nor3_1 _5270_ (.A(_1459_),
    .B(_1461_),
    .C(_1462_),
    .Y(_1463_));
 sky130_fd_sc_hd__or2_1 _5271_ (.A(_1459_),
    .B(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__or2_1 _5272_ (.A(_1434_),
    .B(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__and2_1 _5273_ (.A(_1434_),
    .B(_1464_),
    .X(_1467_));
 sky130_fd_sc_hd__a21oi_1 _5274_ (.A1(_1432_),
    .A2(_1465_),
    .B1(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__xor2_2 _5275_ (.A(_1418_),
    .B(_1468_),
    .X(_1469_));
 sky130_fd_sc_hd__a22o_1 _5276_ (.A1(_0249_),
    .A2(_0671_),
    .B1(_1447_),
    .B2(_1448_),
    .X(_1470_));
 sky130_fd_sc_hd__or3_1 _5277_ (.A(_1437_),
    .B(_1445_),
    .C(_1443_),
    .X(_1471_));
 sky130_fd_sc_hd__o21ai_1 _5278_ (.A1(_1445_),
    .A2(_1443_),
    .B1(_1437_),
    .Y(_1472_));
 sky130_fd_sc_hd__nand2_1 _5279_ (.A(_0726_),
    .B(_0241_),
    .Y(_1473_));
 sky130_fd_sc_hd__and2b_1 _5280_ (.A_N(_1441_),
    .B(_1440_),
    .X(_1474_));
 sky130_fd_sc_hd__xnor2_2 _5281_ (.A(_1473_),
    .B(_1474_),
    .Y(_1475_));
 sky130_fd_sc_hd__and4_1 _5282_ (.A(_0280_),
    .B(_0726_),
    .C(_0531_),
    .D(_0282_),
    .X(_1476_));
 sky130_fd_sc_hd__and2_1 _5283_ (.A(_1475_),
    .B(_1476_),
    .X(_1478_));
 sky130_fd_sc_hd__a21o_1 _5284_ (.A1(_1471_),
    .A2(_1472_),
    .B1(_1478_),
    .X(_1479_));
 sky130_fd_sc_hd__and2_1 _5285_ (.A(_0249_),
    .B(_0506_),
    .X(_1480_));
 sky130_fd_sc_hd__nand3_2 _5286_ (.A(_1471_),
    .B(_1472_),
    .C(_1478_),
    .Y(_1481_));
 sky130_fd_sc_hd__a21bo_1 _5287_ (.A1(_1479_),
    .A2(_1480_),
    .B1_N(_1481_),
    .X(_1482_));
 sky130_fd_sc_hd__nand3_1 _5288_ (.A(_1449_),
    .B(_1470_),
    .C(_1482_),
    .Y(_1483_));
 sky130_fd_sc_hd__and3_1 _5289_ (.A(_1449_),
    .B(_1470_),
    .C(_1482_),
    .X(_1484_));
 sky130_fd_sc_hd__a21oi_1 _5290_ (.A1(_1449_),
    .A2(_1470_),
    .B1(_1482_),
    .Y(_1485_));
 sky130_fd_sc_hd__xnor2_1 _5291_ (.A(_1426_),
    .B(_1428_),
    .Y(_1486_));
 sky130_fd_sc_hd__o2bb2a_1 _5292_ (.A1_N(_0810_),
    .A2_N(_3002_),
    .B1(_1420_),
    .B2(_1421_),
    .X(_1487_));
 sky130_fd_sc_hd__nor2_1 _5293_ (.A(_1423_),
    .B(_1487_),
    .Y(_1489_));
 sky130_fd_sc_hd__and4_1 _5294_ (.A(_0810_),
    .B(_0719_),
    .C(_0293_),
    .D(_0294_),
    .X(_1490_));
 sky130_fd_sc_hd__and2_1 _5295_ (.A(_1489_),
    .B(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__and2_1 _5296_ (.A(_1486_),
    .B(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__nor2_1 _5297_ (.A(_1486_),
    .B(_1491_),
    .Y(_1493_));
 sky130_fd_sc_hd__or2_1 _5298_ (.A(_1492_),
    .B(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__or3_1 _5299_ (.A(_1484_),
    .B(_1485_),
    .C(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__o21a_1 _5300_ (.A1(_1451_),
    .A2(_1454_),
    .B1(_1453_),
    .X(_1496_));
 sky130_fd_sc_hd__a211o_1 _5301_ (.A1(_1483_),
    .A2(_1495_),
    .B1(_1456_),
    .C1(_1496_),
    .X(_1497_));
 sky130_fd_sc_hd__o211ai_2 _5302_ (.A1(_1456_),
    .A2(_1496_),
    .B1(_1483_),
    .C1(_1495_),
    .Y(_1498_));
 sky130_fd_sc_hd__nand3_2 _5303_ (.A(_1492_),
    .B(_1497_),
    .C(_1498_),
    .Y(_1500_));
 sky130_fd_sc_hd__o21a_1 _5304_ (.A1(_1459_),
    .A2(_1462_),
    .B1(_1461_),
    .X(_1501_));
 sky130_fd_sc_hd__a211oi_2 _5305_ (.A1(_1497_),
    .A2(_1500_),
    .B1(_1501_),
    .C1(_1463_),
    .Y(_1502_));
 sky130_fd_sc_hd__xnor2_1 _5306_ (.A(_1434_),
    .B(_1464_),
    .Y(_1503_));
 sky130_fd_sc_hd__xnor2_1 _5307_ (.A(_1432_),
    .B(_1503_),
    .Y(_1504_));
 sky130_fd_sc_hd__o21ai_1 _5308_ (.A1(_1484_),
    .A2(_1485_),
    .B1(_1494_),
    .Y(_1505_));
 sky130_fd_sc_hd__nand3_1 _5309_ (.A(_1481_),
    .B(_1479_),
    .C(_1480_),
    .Y(_1506_));
 sky130_fd_sc_hd__a21o_1 _5310_ (.A1(_1481_),
    .A2(_1479_),
    .B1(_1480_),
    .X(_1507_));
 sky130_fd_sc_hd__xor2_2 _5311_ (.A(_1475_),
    .B(_1476_),
    .X(_1508_));
 sky130_fd_sc_hd__and3_1 _5312_ (.A(_0342_),
    .B(_0421_),
    .C(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__a21o_1 _5313_ (.A1(_1506_),
    .A2(_1507_),
    .B1(_1509_),
    .X(_1511_));
 sky130_fd_sc_hd__nor2_1 _5314_ (.A(_1489_),
    .B(_1490_),
    .Y(_1512_));
 sky130_fd_sc_hd__nor2_1 _5315_ (.A(_1491_),
    .B(_1512_),
    .Y(_1513_));
 sky130_fd_sc_hd__nand3_1 _5316_ (.A(_1506_),
    .B(_1507_),
    .C(_1509_),
    .Y(_1514_));
 sky130_fd_sc_hd__a21bo_1 _5317_ (.A1(_1511_),
    .A2(_1513_),
    .B1_N(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__and3_1 _5318_ (.A(_1495_),
    .B(_1505_),
    .C(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__a21o_1 _5319_ (.A1(_1495_),
    .A2(_1505_),
    .B1(_1515_),
    .X(_1517_));
 sky130_fd_sc_hd__and2b_1 _5320_ (.A_N(_1516_),
    .B(_1517_),
    .X(_1518_));
 sky130_fd_sc_hd__nand3_1 _5321_ (.A(_1514_),
    .B(_1511_),
    .C(_1513_),
    .Y(_1519_));
 sky130_fd_sc_hd__a21o_1 _5322_ (.A1(_1514_),
    .A2(_1511_),
    .B1(_1513_),
    .X(_1520_));
 sky130_fd_sc_hd__nand2_1 _5323_ (.A(_0249_),
    .B(_0421_),
    .Y(_1522_));
 sky130_fd_sc_hd__xnor2_1 _5324_ (.A(_1508_),
    .B(_1522_),
    .Y(_1523_));
 sky130_fd_sc_hd__a22oi_1 _5325_ (.A1(_0280_),
    .A2(_0531_),
    .B1(_0282_),
    .B2(_0964_),
    .Y(_1524_));
 sky130_fd_sc_hd__nor2_1 _5326_ (.A(_1476_),
    .B(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__and3_1 _5327_ (.A(_0342_),
    .B(_0720_),
    .C(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__xnor2_1 _5328_ (.A(_1523_),
    .B(_1526_),
    .Y(_1527_));
 sky130_fd_sc_hd__a22oi_1 _5329_ (.A1(_0720_),
    .A2(_0293_),
    .B1(_0294_),
    .B2(_0810_),
    .Y(_1528_));
 sky130_fd_sc_hd__or2_1 _5330_ (.A(_1490_),
    .B(_1528_),
    .X(_1529_));
 sky130_fd_sc_hd__nor2_1 _5331_ (.A(_1527_),
    .B(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hd__a21o_1 _5332_ (.A1(_1523_),
    .A2(_1526_),
    .B1(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__and3_1 _5333_ (.A(_1519_),
    .B(_1520_),
    .C(_1531_),
    .X(_1533_));
 sky130_fd_sc_hd__a21oi_1 _5334_ (.A1(_1519_),
    .A2(_1520_),
    .B1(_1531_),
    .Y(_1534_));
 sky130_fd_sc_hd__and2_1 _5335_ (.A(_1527_),
    .B(_1529_),
    .X(_1535_));
 sky130_fd_sc_hd__or2_1 _5336_ (.A(_1530_),
    .B(_1535_),
    .X(_1536_));
 sky130_fd_sc_hd__a21oi_1 _5337_ (.A1(_0342_),
    .A2(_0720_),
    .B1(_1525_),
    .Y(_1537_));
 sky130_fd_sc_hd__nor2_1 _5338_ (.A(_1526_),
    .B(_1537_),
    .Y(_1538_));
 sky130_fd_sc_hd__and4_1 _5339_ (.A(_0280_),
    .B(_0964_),
    .C(_0342_),
    .D(_0899_),
    .X(_1539_));
 sky130_fd_sc_hd__nand2_1 _5340_ (.A(_0899_),
    .B(_0293_),
    .Y(_1540_));
 sky130_fd_sc_hd__xnor2_1 _5341_ (.A(_1538_),
    .B(_1539_),
    .Y(_1541_));
 sky130_fd_sc_hd__nor2_1 _5342_ (.A(_1540_),
    .B(_1541_),
    .Y(_1542_));
 sky130_fd_sc_hd__a21oi_1 _5343_ (.A1(_1538_),
    .A2(_1539_),
    .B1(_1542_),
    .Y(_1544_));
 sky130_fd_sc_hd__nor2_1 _5344_ (.A(_1536_),
    .B(_1544_),
    .Y(_1545_));
 sky130_fd_sc_hd__nor3b_1 _5345_ (.A(_1533_),
    .B(_1534_),
    .C_N(_1545_),
    .Y(_1546_));
 sky130_fd_sc_hd__nand2_1 _5346_ (.A(_1518_),
    .B(_1546_),
    .Y(_1547_));
 sky130_fd_sc_hd__a21o_1 _5347_ (.A1(_1497_),
    .A2(_1498_),
    .B1(_1492_),
    .X(_1548_));
 sky130_fd_sc_hd__a21o_1 _5348_ (.A1(_1517_),
    .A2(_1533_),
    .B1(_1516_),
    .X(_1549_));
 sky130_fd_sc_hd__a21oi_1 _5349_ (.A1(_1500_),
    .A2(_1548_),
    .B1(_1549_),
    .Y(_1550_));
 sky130_fd_sc_hd__and3_1 _5350_ (.A(_1500_),
    .B(_1548_),
    .C(_1549_),
    .X(_1551_));
 sky130_fd_sc_hd__nand2_1 _5351_ (.A(_1518_),
    .B(_1533_),
    .Y(_1552_));
 sky130_fd_sc_hd__nand2_1 _5352_ (.A(_1500_),
    .B(_1548_),
    .Y(_1553_));
 sky130_fd_sc_hd__o32ai_4 _5353_ (.A1(_1547_),
    .A2(_1550_),
    .A3(_1551_),
    .B1(_1552_),
    .B2(_1553_),
    .Y(_1555_));
 sky130_fd_sc_hd__o211a_1 _5354_ (.A1(_1463_),
    .A2(_1501_),
    .B1(_1500_),
    .C1(_1497_),
    .X(_1556_));
 sky130_fd_sc_hd__and2_1 _5355_ (.A(_1500_),
    .B(_1548_),
    .X(_1557_));
 sky130_fd_sc_hd__a2bb2o_1 _5356_ (.A1_N(_1502_),
    .A2_N(_1556_),
    .B1(_1557_),
    .B2(_1516_),
    .X(_1558_));
 sky130_fd_sc_hd__and4bb_1 _5357_ (.A_N(_1502_),
    .B_N(_1556_),
    .C(_1557_),
    .D(_1516_),
    .X(_1559_));
 sky130_fd_sc_hd__a21o_1 _5358_ (.A1(_1555_),
    .A2(_1558_),
    .B1(_1559_),
    .X(_1560_));
 sky130_fd_sc_hd__xor2_1 _5359_ (.A(_1504_),
    .B(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__and2_1 _5360_ (.A(_1504_),
    .B(_1560_),
    .X(_1562_));
 sky130_fd_sc_hd__a21oi_2 _5361_ (.A1(_1502_),
    .A2(_1561_),
    .B1(_1562_),
    .Y(_1563_));
 sky130_fd_sc_hd__a21o_1 _5362_ (.A1(_1410_),
    .A2(_1415_),
    .B1(_1350_),
    .X(_1564_));
 sky130_fd_sc_hd__or2b_1 _5363_ (.A(_1468_),
    .B_N(_1418_),
    .X(_1566_));
 sky130_fd_sc_hd__o211ai_4 _5364_ (.A1(_1469_),
    .A2(_1563_),
    .B1(_1564_),
    .C1(_1566_),
    .Y(_1567_));
 sky130_fd_sc_hd__or3b_2 _5365_ (.A(_1349_),
    .B(_1416_),
    .C_N(_1567_),
    .X(_1568_));
 sky130_fd_sc_hd__nand2_1 _5366_ (.A(_1087_),
    .B(_1274_),
    .Y(_1569_));
 sky130_fd_sc_hd__a31o_1 _5367_ (.A1(_1029_),
    .A2(_0506_),
    .A3(_1267_),
    .B1(_1265_),
    .X(_1570_));
 sky130_fd_sc_hd__nor2_1 _5368_ (.A(_1260_),
    .B(_1261_),
    .Y(_1571_));
 sky130_fd_sc_hd__nor2_1 _5369_ (.A(_1262_),
    .B(_1270_),
    .Y(_1572_));
 sky130_fd_sc_hd__nand2_1 _5370_ (.A(_0079_),
    .B(_0671_),
    .Y(_1573_));
 sky130_fd_sc_hd__a31o_1 _5371_ (.A1(_0388_),
    .A2(_0671_),
    .A3(_1247_),
    .B1(_1245_),
    .X(_1574_));
 sky130_fd_sc_hd__and2b_1 _5372_ (.A_N(_1255_),
    .B(_1242_),
    .X(_1575_));
 sky130_fd_sc_hd__nor2_1 _5373_ (.A(_1253_),
    .B(_1575_),
    .Y(_1577_));
 sky130_fd_sc_hd__xnor2_1 _5374_ (.A(_1574_),
    .B(_1577_),
    .Y(_1578_));
 sky130_fd_sc_hd__xnor2_1 _5375_ (.A(_1573_),
    .B(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__a21bo_1 _5376_ (.A1(_1237_),
    .A2(_1239_),
    .B1_N(_1258_),
    .X(_1580_));
 sky130_fd_sc_hd__a21oi_1 _5377_ (.A1(_1249_),
    .A2(_1251_),
    .B1(_1176_),
    .Y(_1581_));
 sky130_fd_sc_hd__and3_1 _5378_ (.A(_1228_),
    .B(_1230_),
    .C(_1232_),
    .X(_1582_));
 sky130_fd_sc_hd__and2b_1 _5379_ (.A_N(_1234_),
    .B(_1153_),
    .X(_1583_));
 sky130_fd_sc_hd__nand2_1 _5380_ (.A(_0388_),
    .B(_0684_),
    .Y(_1584_));
 sky130_fd_sc_hd__buf_2 _5381_ (.A(_0446_),
    .X(_1585_));
 sky130_fd_sc_hd__a21oi_1 _5382_ (.A1(_1585_),
    .A2(_0229_),
    .B1(_1244_),
    .Y(_1586_));
 sky130_fd_sc_hd__and3_1 _5383_ (.A(_1585_),
    .B(_0229_),
    .C(_1244_),
    .X(_1588_));
 sky130_fd_sc_hd__nor2_1 _5384_ (.A(_1586_),
    .B(_1588_),
    .Y(_1589_));
 sky130_fd_sc_hd__xnor2_1 _5385_ (.A(_1584_),
    .B(_1589_),
    .Y(_1590_));
 sky130_fd_sc_hd__o21a_1 _5386_ (.A1(_1582_),
    .A2(_1583_),
    .B1(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__nor3_1 _5387_ (.A(_1582_),
    .B(_1583_),
    .C(_1590_),
    .Y(_1592_));
 sky130_fd_sc_hd__nor2_1 _5388_ (.A(_1591_),
    .B(_1592_),
    .Y(_1593_));
 sky130_fd_sc_hd__xnor2_1 _5389_ (.A(_1581_),
    .B(_1593_),
    .Y(_1594_));
 sky130_fd_sc_hd__and2b_1 _5390_ (.A_N(_1226_),
    .B(_1225_),
    .X(_1595_));
 sky130_fd_sc_hd__clkinv_2 _5391_ (.A(_1236_),
    .Y(_1596_));
 sky130_fd_sc_hd__and2_1 _5392_ (.A(_1227_),
    .B(_1596_),
    .X(_1597_));
 sky130_fd_sc_hd__nand2_2 _5393_ (.A(_0400_),
    .B(_0567_),
    .Y(_1599_));
 sky130_fd_sc_hd__a22o_1 _5394_ (.A1(_0400_),
    .A2(_0697_),
    .B1(_0186_),
    .B2(_0698_),
    .X(_1600_));
 sky130_fd_sc_hd__o21ai_1 _5395_ (.A1(_1220_),
    .A2(_1599_),
    .B1(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__clkbuf_4 _5396_ (.A(_2888_),
    .X(_1602_));
 sky130_fd_sc_hd__a22o_1 _5397_ (.A1(_1602_),
    .A2(_0573_),
    .B1(_0581_),
    .B2(_1229_),
    .X(_1603_));
 sky130_fd_sc_hd__nand2_1 _5398_ (.A(_0573_),
    .B(_1231_),
    .Y(_1604_));
 sky130_fd_sc_hd__nand2_1 _5399_ (.A(_1603_),
    .B(_1604_),
    .Y(_1605_));
 sky130_fd_sc_hd__a31o_1 _5400_ (.A1(_0400_),
    .A2(_0573_),
    .A3(_1222_),
    .B1(_1221_),
    .X(_1606_));
 sky130_fd_sc_hd__xor2_1 _5401_ (.A(_1605_),
    .B(_1606_),
    .X(_1607_));
 sky130_fd_sc_hd__xor2_1 _5402_ (.A(_1232_),
    .B(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__xnor2_1 _5403_ (.A(_1601_),
    .B(_1608_),
    .Y(_1610_));
 sky130_fd_sc_hd__o21ai_1 _5404_ (.A1(_1595_),
    .A2(_1597_),
    .B1(_1610_),
    .Y(_1611_));
 sky130_fd_sc_hd__or3_1 _5405_ (.A(_1595_),
    .B(_1597_),
    .C(_1610_),
    .X(_1612_));
 sky130_fd_sc_hd__and2_1 _5406_ (.A(_1611_),
    .B(_1612_),
    .X(_1613_));
 sky130_fd_sc_hd__xnor2_1 _5407_ (.A(_1594_),
    .B(_1613_),
    .Y(_1614_));
 sky130_fd_sc_hd__xor2_1 _5408_ (.A(_1580_),
    .B(_1614_),
    .X(_1615_));
 sky130_fd_sc_hd__xnor2_1 _5409_ (.A(_1579_),
    .B(_1615_),
    .Y(_1616_));
 sky130_fd_sc_hd__o21ai_1 _5410_ (.A1(_1571_),
    .A2(_1572_),
    .B1(_1616_),
    .Y(_1617_));
 sky130_fd_sc_hd__or3_1 _5411_ (.A(_1571_),
    .B(_1572_),
    .C(_1616_),
    .X(_1618_));
 sky130_fd_sc_hd__and2_1 _5412_ (.A(_1617_),
    .B(_1618_),
    .X(_1619_));
 sky130_fd_sc_hd__xnor2_1 _5413_ (.A(_1570_),
    .B(_1619_),
    .Y(_1621_));
 sky130_fd_sc_hd__a21oi_1 _5414_ (.A1(_1272_),
    .A2(_1569_),
    .B1(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__and3_1 _5415_ (.A(_1272_),
    .B(_1569_),
    .C(_1621_),
    .X(_1623_));
 sky130_fd_sc_hd__nor2_1 _5416_ (.A(_1622_),
    .B(_1623_),
    .Y(_1624_));
 sky130_fd_sc_hd__a21oi_1 _5417_ (.A1(_1348_),
    .A2(_1568_),
    .B1(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__or2_1 _5418_ (.A(net15),
    .B(_2883_),
    .X(_1626_));
 sky130_fd_sc_hd__clkbuf_4 _5419_ (.A(_1626_),
    .X(_1627_));
 sky130_fd_sc_hd__a31o_1 _5420_ (.A1(_1348_),
    .A2(_1568_),
    .A3(_1624_),
    .B1(_1627_),
    .X(_1628_));
 sky130_fd_sc_hd__or2_2 _5421_ (.A(_1625_),
    .B(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__o211a_1 _5422_ (.A1(_2881_),
    .A2(_1027_),
    .B1(_1028_),
    .C1(_1629_),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 _5423_ (.A(_1627_),
    .X(_1631_));
 sky130_fd_sc_hd__a21o_1 _5424_ (.A1(_1272_),
    .A2(_1569_),
    .B1(_1621_),
    .X(_1632_));
 sky130_fd_sc_hd__nand2_1 _5425_ (.A(_1570_),
    .B(_1619_),
    .Y(_1633_));
 sky130_fd_sc_hd__nand2_1 _5426_ (.A(_1594_),
    .B(_1613_),
    .Y(_1634_));
 sky130_fd_sc_hd__and2b_1 _5427_ (.A_N(_1601_),
    .B(_1608_),
    .X(_1635_));
 sky130_fd_sc_hd__nor2_1 _5428_ (.A(_1220_),
    .B(_1599_),
    .Y(_1636_));
 sky130_fd_sc_hd__nand2_1 _5429_ (.A(_1229_),
    .B(_0572_),
    .Y(_1637_));
 sky130_fd_sc_hd__nand2_1 _5430_ (.A(_2888_),
    .B(_0568_),
    .Y(_1638_));
 sky130_fd_sc_hd__xor2_1 _5431_ (.A(_1637_),
    .B(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__xnor2_1 _5432_ (.A(_1636_),
    .B(_1639_),
    .Y(_1640_));
 sky130_fd_sc_hd__and2_1 _5433_ (.A(_1604_),
    .B(_1640_),
    .X(_1642_));
 sky130_fd_sc_hd__nor2_1 _5434_ (.A(_1604_),
    .B(_1640_),
    .Y(_1643_));
 sky130_fd_sc_hd__or2_1 _5435_ (.A(_1642_),
    .B(_1643_),
    .X(_1644_));
 sky130_fd_sc_hd__xor2_1 _5436_ (.A(_1599_),
    .B(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__or2_1 _5437_ (.A(_1635_),
    .B(_1645_),
    .X(_1646_));
 sky130_fd_sc_hd__nand2_1 _5438_ (.A(_1635_),
    .B(_1645_),
    .Y(_1647_));
 sky130_fd_sc_hd__nand2_1 _5439_ (.A(_1646_),
    .B(_1647_),
    .Y(_1648_));
 sky130_fd_sc_hd__nor2_1 _5440_ (.A(_1232_),
    .B(_1607_),
    .Y(_1649_));
 sky130_fd_sc_hd__a31o_1 _5441_ (.A1(_1603_),
    .A2(_1604_),
    .A3(_1606_),
    .B1(_1649_),
    .X(_1650_));
 sky130_fd_sc_hd__a22o_1 _5442_ (.A1(_0378_),
    .A2(_1585_),
    .B1(_0388_),
    .B2(_0546_),
    .X(_1651_));
 sky130_fd_sc_hd__inv_2 _5443_ (.A(_1651_),
    .Y(_1653_));
 sky130_fd_sc_hd__and3_1 _5444_ (.A(_1585_),
    .B(_0388_),
    .C(_1244_),
    .X(_1654_));
 sky130_fd_sc_hd__nor2_1 _5445_ (.A(_1653_),
    .B(_1654_),
    .Y(_1655_));
 sky130_fd_sc_hd__xnor2_1 _5446_ (.A(_1650_),
    .B(_1655_),
    .Y(_1656_));
 sky130_fd_sc_hd__or2_1 _5447_ (.A(_1648_),
    .B(_1656_),
    .X(_1657_));
 sky130_fd_sc_hd__nand2_1 _5448_ (.A(_1648_),
    .B(_1656_),
    .Y(_1658_));
 sky130_fd_sc_hd__nand2_1 _5449_ (.A(_1657_),
    .B(_1658_),
    .Y(_1659_));
 sky130_fd_sc_hd__a21o_1 _5450_ (.A1(_1611_),
    .A2(_1634_),
    .B1(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__nand3_1 _5451_ (.A(_1611_),
    .B(_1634_),
    .C(_1659_),
    .Y(_1661_));
 sky130_fd_sc_hd__and2_1 _5452_ (.A(_1660_),
    .B(_1661_),
    .X(_1662_));
 sky130_fd_sc_hd__and2b_1 _5453_ (.A_N(_1581_),
    .B(_1593_),
    .X(_1664_));
 sky130_fd_sc_hd__o21ba_1 _5454_ (.A1(_1584_),
    .A2(_1586_),
    .B1_N(_1588_),
    .X(_1665_));
 sky130_fd_sc_hd__o21ba_1 _5455_ (.A1(_1591_),
    .A2(_1664_),
    .B1_N(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__or3b_1 _5456_ (.A(_1591_),
    .B(_1664_),
    .C_N(_1665_),
    .X(_1667_));
 sky130_fd_sc_hd__and2b_1 _5457_ (.A_N(_1666_),
    .B(_1667_),
    .X(_1668_));
 sky130_fd_sc_hd__nand2_1 _5458_ (.A(_0079_),
    .B(_0684_),
    .Y(_1669_));
 sky130_fd_sc_hd__xnor2_1 _5459_ (.A(_1668_),
    .B(_1669_),
    .Y(_1670_));
 sky130_fd_sc_hd__xnor2_1 _5460_ (.A(_1662_),
    .B(_1670_),
    .Y(_1671_));
 sky130_fd_sc_hd__or2b_1 _5461_ (.A(_1580_),
    .B_N(_1614_),
    .X(_1672_));
 sky130_fd_sc_hd__and2b_1 _5462_ (.A_N(_1614_),
    .B(_1580_),
    .X(_1673_));
 sky130_fd_sc_hd__a21o_1 _5463_ (.A1(_1579_),
    .A2(_1672_),
    .B1(_1673_),
    .X(_1675_));
 sky130_fd_sc_hd__xor2_1 _5464_ (.A(_1671_),
    .B(_1675_),
    .X(_1676_));
 sky130_fd_sc_hd__o21ai_1 _5465_ (.A1(_1253_),
    .A2(_1575_),
    .B1(_1574_),
    .Y(_1677_));
 sky130_fd_sc_hd__or2b_1 _5466_ (.A(_1573_),
    .B_N(_1578_),
    .X(_1678_));
 sky130_fd_sc_hd__nand2_1 _5467_ (.A(_1677_),
    .B(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__xor2_1 _5468_ (.A(_1676_),
    .B(_1679_),
    .X(_1680_));
 sky130_fd_sc_hd__a21oi_1 _5469_ (.A1(_1617_),
    .A2(_1633_),
    .B1(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__and3_1 _5470_ (.A(_1617_),
    .B(_1633_),
    .C(_1680_),
    .X(_1682_));
 sky130_fd_sc_hd__or2_1 _5471_ (.A(_1681_),
    .B(_1682_),
    .X(_1683_));
 sky130_fd_sc_hd__a311oi_4 _5472_ (.A1(_1348_),
    .A2(_1568_),
    .A3(_1632_),
    .B1(_1623_),
    .C1(_1683_),
    .Y(_1684_));
 sky130_fd_sc_hd__a31o_1 _5473_ (.A1(_1348_),
    .A2(_1568_),
    .A3(_1632_),
    .B1(_1623_),
    .X(_1686_));
 sky130_fd_sc_hd__and2_1 _5474_ (.A(_1683_),
    .B(_1686_),
    .X(_1687_));
 sky130_fd_sc_hd__nor2_2 _5475_ (.A(_1684_),
    .B(_1687_),
    .Y(_1688_));
 sky130_fd_sc_hd__and3_1 _5476_ (.A(_0696_),
    .B(_0671_),
    .C(_0678_),
    .X(_1689_));
 sky130_fd_sc_hd__a21oi_2 _5477_ (.A1(_0675_),
    .A2(_0677_),
    .B1(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hd__and2b_1 _5478_ (.A_N(_0712_),
    .B(_0681_),
    .X(_1691_));
 sky130_fd_sc_hd__and2b_1 _5479_ (.A_N(_0679_),
    .B(_0713_),
    .X(_1692_));
 sky130_fd_sc_hd__and3_1 _5480_ (.A(_0699_),
    .B(_0700_),
    .C(_0709_),
    .X(_1693_));
 sky130_fd_sc_hd__nand2_1 _5481_ (.A(_0567_),
    .B(_2856_),
    .Y(_1694_));
 sky130_fd_sc_hd__nand2_1 _5482_ (.A(_0568_),
    .B(_0740_),
    .Y(_1695_));
 sky130_fd_sc_hd__xor2_1 _5483_ (.A(_0703_),
    .B(_1695_),
    .X(_1697_));
 sky130_fd_sc_hd__xor2_1 _5484_ (.A(_0700_),
    .B(_1697_),
    .X(_1698_));
 sky130_fd_sc_hd__xnor2_1 _5485_ (.A(_0704_),
    .B(_1698_),
    .Y(_1699_));
 sky130_fd_sc_hd__or2_1 _5486_ (.A(_1694_),
    .B(_1699_),
    .X(_1700_));
 sky130_fd_sc_hd__nand2_1 _5487_ (.A(_1694_),
    .B(_1699_),
    .Y(_1701_));
 sky130_fd_sc_hd__and2_1 _5488_ (.A(_1700_),
    .B(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__xnor2_1 _5489_ (.A(_1693_),
    .B(_1702_),
    .Y(_1703_));
 sky130_fd_sc_hd__inv_2 _5490_ (.A(_0583_),
    .Y(_1704_));
 sky130_fd_sc_hd__nor2_1 _5491_ (.A(_1704_),
    .B(_0708_),
    .Y(_1705_));
 sky130_fd_sc_hd__a31o_1 _5492_ (.A1(_0702_),
    .A2(_0704_),
    .A3(_0706_),
    .B1(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__nand2_1 _5493_ (.A(_1585_),
    .B(_2833_),
    .Y(_1708_));
 sky130_fd_sc_hd__a22o_1 _5494_ (.A1(_1585_),
    .A2(_1521_),
    .B1(_2833_),
    .B2(_0546_),
    .X(_1709_));
 sky130_fd_sc_hd__o21a_1 _5495_ (.A1(_0545_),
    .A2(_1708_),
    .B1(_1709_),
    .X(_1710_));
 sky130_fd_sc_hd__xnor2_1 _5496_ (.A(_1706_),
    .B(_1710_),
    .Y(_1711_));
 sky130_fd_sc_hd__or2_1 _5497_ (.A(_1703_),
    .B(_1711_),
    .X(_1712_));
 sky130_fd_sc_hd__nand2_1 _5498_ (.A(_1703_),
    .B(_1711_),
    .Y(_1713_));
 sky130_fd_sc_hd__nand2_1 _5499_ (.A(_1712_),
    .B(_1713_),
    .Y(_1714_));
 sky130_fd_sc_hd__or2b_1 _5500_ (.A(_0695_),
    .B_N(_0710_),
    .X(_1715_));
 sky130_fd_sc_hd__a21bo_1 _5501_ (.A1(_0694_),
    .A2(_0711_),
    .B1_N(_1715_),
    .X(_1716_));
 sky130_fd_sc_hd__xor2_1 _5502_ (.A(_1714_),
    .B(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__and2b_1 _5503_ (.A_N(_0682_),
    .B(_0693_),
    .X(_1719_));
 sky130_fd_sc_hd__o21ba_1 _5504_ (.A1(_0686_),
    .A2(_0687_),
    .B1_N(_0688_),
    .X(_1720_));
 sky130_fd_sc_hd__o21ba_1 _5505_ (.A1(_0691_),
    .A2(_1719_),
    .B1_N(_1720_),
    .X(_1721_));
 sky130_fd_sc_hd__or3b_1 _5506_ (.A(_0691_),
    .B(_1719_),
    .C_N(_1720_),
    .X(_1722_));
 sky130_fd_sc_hd__and2b_1 _5507_ (.A_N(_1721_),
    .B(_1722_),
    .X(_1723_));
 sky130_fd_sc_hd__nand2_1 _5508_ (.A(_0684_),
    .B(_0674_),
    .Y(_1724_));
 sky130_fd_sc_hd__xor2_1 _5509_ (.A(_1723_),
    .B(_1724_),
    .X(_1725_));
 sky130_fd_sc_hd__xor2_1 _5510_ (.A(_1717_),
    .B(_1725_),
    .X(_1726_));
 sky130_fd_sc_hd__o21ai_2 _5511_ (.A1(_1691_),
    .A2(_1692_),
    .B1(_1726_),
    .Y(_1727_));
 sky130_fd_sc_hd__or3_1 _5512_ (.A(_1691_),
    .B(_1692_),
    .C(_1726_),
    .X(_1728_));
 sky130_fd_sc_hd__and2_1 _5513_ (.A(_1727_),
    .B(_1728_),
    .X(_1730_));
 sky130_fd_sc_hd__xnor2_2 _5514_ (.A(_1690_),
    .B(_1730_),
    .Y(_1731_));
 sky130_fd_sc_hd__and2b_1 _5515_ (.A_N(_0668_),
    .B(_0715_),
    .X(_1732_));
 sky130_fd_sc_hd__o21ba_1 _5516_ (.A1(_0670_),
    .A2(_0714_),
    .B1_N(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__xor2_2 _5517_ (.A(_1731_),
    .B(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__nand3b_1 _5518_ (.A_N(_0717_),
    .B(_1020_),
    .C(_1019_),
    .Y(_1735_));
 sky130_fd_sc_hd__or4b_1 _5519_ (.A(_0717_),
    .B(_1000_),
    .C(_1013_),
    .D_N(_1020_),
    .X(_1736_));
 sky130_fd_sc_hd__a22o_1 _5520_ (.A1(_0667_),
    .A2(_0716_),
    .B1(_0796_),
    .B2(_0797_),
    .X(_1737_));
 sky130_fd_sc_hd__o21a_1 _5521_ (.A1(_0667_),
    .A2(_0716_),
    .B1(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__inv_2 _5522_ (.A(_1738_),
    .Y(_1739_));
 sky130_fd_sc_hd__nand4_1 _5523_ (.A(_1734_),
    .B(_1735_),
    .C(_1736_),
    .D(_1739_),
    .Y(_1741_));
 sky130_fd_sc_hd__a31o_2 _5524_ (.A1(_1735_),
    .A2(_1736_),
    .A3(_1739_),
    .B1(_1734_),
    .X(_1742_));
 sky130_fd_sc_hd__and2_1 _5525_ (.A(_2882_),
    .B(_2883_),
    .X(_1743_));
 sky130_fd_sc_hd__clkbuf_2 _5526_ (.A(_1743_),
    .X(_1744_));
 sky130_fd_sc_hd__and3_1 _5527_ (.A(_1741_),
    .B(_1742_),
    .C(_1744_),
    .X(_1745_));
 sky130_fd_sc_hd__and2b_1 _5528_ (.A_N(_0414_),
    .B(_0376_),
    .X(_1746_));
 sky130_fd_sc_hd__and2_1 _5529_ (.A(_0374_),
    .B(_0415_),
    .X(_1747_));
 sky130_fd_sc_hd__o21ba_1 _5530_ (.A1(_0379_),
    .A2(_2999_),
    .B1_N(_0381_),
    .X(_1748_));
 sky130_fd_sc_hd__a31o_1 _5531_ (.A1(_1029_),
    .A2(_2668_),
    .A3(_0382_),
    .B1(_1748_),
    .X(_1749_));
 sky130_fd_sc_hd__and2b_1 _5532_ (.A_N(_0402_),
    .B(_0409_),
    .X(_1750_));
 sky130_fd_sc_hd__nor2_1 _5533_ (.A(_3021_),
    .B(_0399_),
    .Y(_1752_));
 sky130_fd_sc_hd__nand2_1 _5534_ (.A(_2888_),
    .B(_2858_),
    .Y(_1753_));
 sky130_fd_sc_hd__xor2_1 _5535_ (.A(_0404_),
    .B(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__xnor2_1 _5536_ (.A(_1752_),
    .B(_1754_),
    .Y(_1755_));
 sky130_fd_sc_hd__and2_1 _5537_ (.A(_0405_),
    .B(_1755_),
    .X(_1756_));
 sky130_fd_sc_hd__nor2_1 _5538_ (.A(_0405_),
    .B(_1755_),
    .Y(_1757_));
 sky130_fd_sc_hd__or2_1 _5539_ (.A(_1756_),
    .B(_1757_),
    .X(_1758_));
 sky130_fd_sc_hd__xor2_1 _5540_ (.A(_0399_),
    .B(_1758_),
    .X(_1759_));
 sky130_fd_sc_hd__xnor2_1 _5541_ (.A(_1750_),
    .B(_1759_),
    .Y(_1760_));
 sky130_fd_sc_hd__inv_2 _5542_ (.A(_3032_),
    .Y(_1761_));
 sky130_fd_sc_hd__nor2_1 _5543_ (.A(_1761_),
    .B(_0408_),
    .Y(_1763_));
 sky130_fd_sc_hd__a31o_1 _5544_ (.A1(_0403_),
    .A2(_0405_),
    .A3(_0407_),
    .B1(_1763_),
    .X(_1764_));
 sky130_fd_sc_hd__a22o_1 _5545_ (.A1(_0378_),
    .A2(_2845_),
    .B1(_2551_),
    .B2(_0388_),
    .X(_1765_));
 sky130_fd_sc_hd__inv_2 _5546_ (.A(_1765_),
    .Y(_1766_));
 sky130_fd_sc_hd__and4_1 _5547_ (.A(_0378_),
    .B(_0388_),
    .C(_2845_),
    .D(_2551_),
    .X(_1767_));
 sky130_fd_sc_hd__nor2_1 _5548_ (.A(_1766_),
    .B(_1767_),
    .Y(_1768_));
 sky130_fd_sc_hd__xnor2_1 _5549_ (.A(_1764_),
    .B(_1768_),
    .Y(_1769_));
 sky130_fd_sc_hd__or2_1 _5550_ (.A(_1760_),
    .B(_1769_),
    .X(_1770_));
 sky130_fd_sc_hd__nand2_1 _5551_ (.A(_1760_),
    .B(_1769_),
    .Y(_1771_));
 sky130_fd_sc_hd__nand2_1 _5552_ (.A(_1770_),
    .B(_1771_),
    .Y(_1772_));
 sky130_fd_sc_hd__or2b_1 _5553_ (.A(_0398_),
    .B_N(_0410_),
    .X(_1774_));
 sky130_fd_sc_hd__a21bo_1 _5554_ (.A1(_0397_),
    .A2(_0411_),
    .B1_N(_1774_),
    .X(_1775_));
 sky130_fd_sc_hd__xnor2_1 _5555_ (.A(_1772_),
    .B(_1775_),
    .Y(_1776_));
 sky130_fd_sc_hd__and2b_1 _5556_ (.A_N(_0386_),
    .B(_0396_),
    .X(_1777_));
 sky130_fd_sc_hd__o21ba_1 _5557_ (.A1(_0389_),
    .A2(_0390_),
    .B1_N(_0391_),
    .X(_1778_));
 sky130_fd_sc_hd__o21ba_1 _5558_ (.A1(_0394_),
    .A2(_1777_),
    .B1_N(_1778_),
    .X(_1779_));
 sky130_fd_sc_hd__or3b_1 _5559_ (.A(_0394_),
    .B(_1777_),
    .C_N(_1778_),
    .X(_1780_));
 sky130_fd_sc_hd__and2b_1 _5560_ (.A_N(_1779_),
    .B(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__nand2_1 _5561_ (.A(_2886_),
    .B(_2676_),
    .Y(_1782_));
 sky130_fd_sc_hd__xnor2_1 _5562_ (.A(_1781_),
    .B(_1782_),
    .Y(_1783_));
 sky130_fd_sc_hd__xnor2_1 _5563_ (.A(_1776_),
    .B(_1783_),
    .Y(_1785_));
 sky130_fd_sc_hd__nor2_1 _5564_ (.A(_0385_),
    .B(_0412_),
    .Y(_1786_));
 sky130_fd_sc_hd__a21o_1 _5565_ (.A1(_0383_),
    .A2(_0413_),
    .B1(_1786_),
    .X(_1787_));
 sky130_fd_sc_hd__xor2_1 _5566_ (.A(_1785_),
    .B(_1787_),
    .X(_1788_));
 sky130_fd_sc_hd__xnor2_1 _5567_ (.A(_1749_),
    .B(_1788_),
    .Y(_1789_));
 sky130_fd_sc_hd__o21ai_1 _5568_ (.A1(_1746_),
    .A2(_1747_),
    .B1(_1789_),
    .Y(_1790_));
 sky130_fd_sc_hd__or3_1 _5569_ (.A(_1746_),
    .B(_1747_),
    .C(_1789_),
    .X(_1791_));
 sky130_fd_sc_hd__nand2_1 _5570_ (.A(_1790_),
    .B(_1791_),
    .Y(_1792_));
 sky130_fd_sc_hd__or2_1 _5571_ (.A(_0149_),
    .B(_0417_),
    .X(_1793_));
 sky130_fd_sc_hd__a211o_1 _5572_ (.A1(_0368_),
    .A2(_0366_),
    .B1(_1793_),
    .C1(_0218_),
    .X(_1794_));
 sky130_fd_sc_hd__or2b_1 _5573_ (.A(_0218_),
    .B_N(_0368_),
    .X(_1796_));
 sky130_fd_sc_hd__or4_1 _5574_ (.A(_0361_),
    .B(_0365_),
    .C(_1796_),
    .D(_1793_),
    .X(_1797_));
 sky130_fd_sc_hd__o22a_1 _5575_ (.A1(_0078_),
    .A2(_0148_),
    .B1(_0373_),
    .B2(_0416_),
    .X(_1798_));
 sky130_fd_sc_hd__a21o_1 _5576_ (.A1(_0373_),
    .A2(_0416_),
    .B1(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__and4_1 _5577_ (.A(_1792_),
    .B(_1794_),
    .C(_1797_),
    .D(_1799_),
    .X(_1800_));
 sky130_fd_sc_hd__a31o_1 _5578_ (.A1(_1794_),
    .A2(_1797_),
    .A3(_1799_),
    .B1(_1792_),
    .X(_1801_));
 sky130_fd_sc_hd__nand2_1 _5579_ (.A(_2885_),
    .B(_1801_),
    .Y(_1802_));
 sky130_fd_sc_hd__and2b_1 _5580_ (.A_N(_2874_),
    .B(_2832_),
    .X(_1803_));
 sky130_fd_sc_hd__and2_1 _5581_ (.A(_2830_),
    .B(_2875_),
    .X(_1804_));
 sky130_fd_sc_hd__a21o_1 _5582_ (.A1(_2834_),
    .A2(_2835_),
    .B1(_2837_),
    .X(_1805_));
 sky130_fd_sc_hd__and2b_1 _5583_ (.A_N(_2861_),
    .B(_2869_),
    .X(_1807_));
 sky130_fd_sc_hd__nor2_1 _5584_ (.A(_2442_),
    .B(_2857_),
    .Y(_1808_));
 sky130_fd_sc_hd__nand2_1 _5585_ (.A(_2405_),
    .B(_0740_),
    .Y(_1809_));
 sky130_fd_sc_hd__xor2_1 _5586_ (.A(_2864_),
    .B(_1809_),
    .X(_1810_));
 sky130_fd_sc_hd__xnor2_1 _5587_ (.A(_1808_),
    .B(_1810_),
    .Y(_1811_));
 sky130_fd_sc_hd__and2_1 _5588_ (.A(_2865_),
    .B(_1811_),
    .X(_1812_));
 sky130_fd_sc_hd__nor2_1 _5589_ (.A(_2865_),
    .B(_1811_),
    .Y(_1813_));
 sky130_fd_sc_hd__or2_1 _5590_ (.A(_1812_),
    .B(_1813_),
    .X(_1814_));
 sky130_fd_sc_hd__xor2_1 _5591_ (.A(_2857_),
    .B(_1814_),
    .X(_1815_));
 sky130_fd_sc_hd__xnor2_1 _5592_ (.A(_1807_),
    .B(_1815_),
    .Y(_1816_));
 sky130_fd_sc_hd__inv_2 _5593_ (.A(_2454_),
    .Y(_1818_));
 sky130_fd_sc_hd__nor2_1 _5594_ (.A(_1818_),
    .B(_2868_),
    .Y(_1819_));
 sky130_fd_sc_hd__a31o_1 _5595_ (.A1(_2863_),
    .A2(_2865_),
    .A3(_2867_),
    .B1(_1819_),
    .X(_1820_));
 sky130_fd_sc_hd__a22o_1 _5596_ (.A1(_2845_),
    .A2(_1521_),
    .B1(_2551_),
    .B2(_2833_),
    .X(_1821_));
 sky130_fd_sc_hd__inv_2 _5597_ (.A(_1821_),
    .Y(_1822_));
 sky130_fd_sc_hd__and3_1 _5598_ (.A(_2845_),
    .B(_2833_),
    .C(_2846_),
    .X(_1823_));
 sky130_fd_sc_hd__nor2_1 _5599_ (.A(_1822_),
    .B(_1823_),
    .Y(_1824_));
 sky130_fd_sc_hd__xnor2_1 _5600_ (.A(_1820_),
    .B(_1824_),
    .Y(_1825_));
 sky130_fd_sc_hd__or2_1 _5601_ (.A(_1816_),
    .B(_1825_),
    .X(_1826_));
 sky130_fd_sc_hd__nand2_1 _5602_ (.A(_1816_),
    .B(_1825_),
    .Y(_1827_));
 sky130_fd_sc_hd__nand2_1 _5603_ (.A(_1826_),
    .B(_1827_),
    .Y(_1829_));
 sky130_fd_sc_hd__or2b_1 _5604_ (.A(_2855_),
    .B_N(_2870_),
    .X(_1830_));
 sky130_fd_sc_hd__a21bo_1 _5605_ (.A1(_2854_),
    .A2(_2871_),
    .B1_N(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__xnor2_1 _5606_ (.A(_1829_),
    .B(_1831_),
    .Y(_1832_));
 sky130_fd_sc_hd__and2b_1 _5607_ (.A_N(_2842_),
    .B(_2853_),
    .X(_1833_));
 sky130_fd_sc_hd__o21ba_1 _5608_ (.A1(_2844_),
    .A2(_2847_),
    .B1_N(_2848_),
    .X(_1834_));
 sky130_fd_sc_hd__o21ba_1 _5609_ (.A1(_2851_),
    .A2(_1833_),
    .B1_N(_1834_),
    .X(_1835_));
 sky130_fd_sc_hd__or3b_1 _5610_ (.A(_2851_),
    .B(_1833_),
    .C_N(_1834_),
    .X(_1836_));
 sky130_fd_sc_hd__and2b_1 _5611_ (.A_N(_1835_),
    .B(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__nand2_1 _5612_ (.A(_2676_),
    .B(_0674_),
    .Y(_1838_));
 sky130_fd_sc_hd__xnor2_1 _5613_ (.A(_1837_),
    .B(_1838_),
    .Y(_1840_));
 sky130_fd_sc_hd__xnor2_1 _5614_ (.A(_1832_),
    .B(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__nor2_1 _5615_ (.A(_2841_),
    .B(_2872_),
    .Y(_1842_));
 sky130_fd_sc_hd__a21o_1 _5616_ (.A1(_2839_),
    .A2(_2873_),
    .B1(_1842_),
    .X(_1843_));
 sky130_fd_sc_hd__xor2_1 _5617_ (.A(_1841_),
    .B(_1843_),
    .X(_1844_));
 sky130_fd_sc_hd__xnor2_2 _5618_ (.A(_1805_),
    .B(_1844_),
    .Y(_1845_));
 sky130_fd_sc_hd__o21ai_2 _5619_ (.A1(_1803_),
    .A2(_1804_),
    .B1(_1845_),
    .Y(_1846_));
 sky130_fd_sc_hd__or3_1 _5620_ (.A(_1803_),
    .B(_1804_),
    .C(_1845_),
    .X(_1847_));
 sky130_fd_sc_hd__nand2_1 _5621_ (.A(_1846_),
    .B(_1847_),
    .Y(_1848_));
 sky130_fd_sc_hd__nand2_1 _5622_ (.A(_2617_),
    .B(_2877_),
    .Y(_1849_));
 sky130_fd_sc_hd__or2b_1 _5623_ (.A(_1849_),
    .B_N(_2824_),
    .X(_1851_));
 sky130_fd_sc_hd__nand2_1 _5624_ (.A(_2818_),
    .B(_2822_),
    .Y(_1852_));
 sky130_fd_sc_hd__or3b_1 _5625_ (.A(_1852_),
    .B(_1849_),
    .C_N(_2811_),
    .X(_1853_));
 sky130_fd_sc_hd__a21o_1 _5626_ (.A1(_2829_),
    .A2(_2876_),
    .B1(_2826_),
    .X(_1854_));
 sky130_fd_sc_hd__o21a_1 _5627_ (.A1(_2829_),
    .A2(_2876_),
    .B1(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__a31o_2 _5628_ (.A1(_1851_),
    .A2(_1853_),
    .A3(_1855_),
    .B1(_1848_),
    .X(_1856_));
 sky130_fd_sc_hd__nand2_1 _5629_ (.A(_2879_),
    .B(_1856_),
    .Y(_1857_));
 sky130_fd_sc_hd__a41o_1 _5630_ (.A1(_1848_),
    .A2(_1851_),
    .A3(_1853_),
    .A4(_1855_),
    .B1(_1857_),
    .X(_1858_));
 sky130_fd_sc_hd__o21ai_1 _5631_ (.A1(_1800_),
    .A2(_1802_),
    .B1(_1858_),
    .Y(_1859_));
 sky130_fd_sc_hd__or3_1 _5632_ (.A(_1024_),
    .B(_1745_),
    .C(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__clkbuf_4 _5633_ (.A(_1028_),
    .X(_1862_));
 sky130_fd_sc_hd__o211a_1 _5634_ (.A1(_1631_),
    .A2(_1688_),
    .B1(_1860_),
    .C1(_1862_),
    .X(net19));
 sky130_fd_sc_hd__and2b_1 _5635_ (.A_N(_1671_),
    .B(_1675_),
    .X(_1863_));
 sky130_fd_sc_hd__and2b_1 _5636_ (.A_N(_1676_),
    .B(_1679_),
    .X(_1864_));
 sky130_fd_sc_hd__nand2_1 _5637_ (.A(_1662_),
    .B(_1670_),
    .Y(_1865_));
 sky130_fd_sc_hd__nand2_1 _5638_ (.A(_0698_),
    .B(_1602_),
    .Y(_1866_));
 sky130_fd_sc_hd__nand2_1 _5639_ (.A(_1602_),
    .B(_0573_),
    .Y(_1867_));
 sky130_fd_sc_hd__and3_1 _5640_ (.A(_0697_),
    .B(_1229_),
    .C(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__xor2_1 _5641_ (.A(_1866_),
    .B(_1868_),
    .X(_1869_));
 sky130_fd_sc_hd__o21a_1 _5642_ (.A1(_1599_),
    .A2(_1644_),
    .B1(_1869_),
    .X(_1870_));
 sky130_fd_sc_hd__nor3_1 _5643_ (.A(_1599_),
    .B(_1644_),
    .C(_1869_),
    .Y(_1872_));
 sky130_fd_sc_hd__or2_1 _5644_ (.A(_1870_),
    .B(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__nand2_1 _5645_ (.A(_1585_),
    .B(_0388_),
    .Y(_1874_));
 sky130_fd_sc_hd__a21oi_1 _5646_ (.A1(_1636_),
    .A2(_1639_),
    .B1(_1643_),
    .Y(_1875_));
 sky130_fd_sc_hd__xnor2_1 _5647_ (.A(_1874_),
    .B(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__nor2_1 _5648_ (.A(_1873_),
    .B(_1876_),
    .Y(_1877_));
 sky130_fd_sc_hd__and2_1 _5649_ (.A(_1873_),
    .B(_1876_),
    .X(_1878_));
 sky130_fd_sc_hd__or2_1 _5650_ (.A(_1877_),
    .B(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__a21oi_1 _5651_ (.A1(_1647_),
    .A2(_1657_),
    .B1(_1879_),
    .Y(_1880_));
 sky130_fd_sc_hd__and3_1 _5652_ (.A(_1647_),
    .B(_1657_),
    .C(_1879_),
    .X(_1881_));
 sky130_fd_sc_hd__or2_1 _5653_ (.A(_1880_),
    .B(_1881_),
    .X(_1883_));
 sky130_fd_sc_hd__o21ai_1 _5654_ (.A1(_1650_),
    .A2(_1654_),
    .B1(_1651_),
    .Y(_1884_));
 sky130_fd_sc_hd__and3b_1 _5655_ (.A_N(_1884_),
    .B(_0079_),
    .C(_0546_),
    .X(_1885_));
 sky130_fd_sc_hd__a21bo_1 _5656_ (.A1(_0546_),
    .A2(_0079_),
    .B1_N(_1884_),
    .X(_1886_));
 sky130_fd_sc_hd__or2b_1 _5657_ (.A(_1885_),
    .B_N(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__nor2_1 _5658_ (.A(_1883_),
    .B(_1887_),
    .Y(_1888_));
 sky130_fd_sc_hd__and2_1 _5659_ (.A(_1883_),
    .B(_1887_),
    .X(_1889_));
 sky130_fd_sc_hd__or2_1 _5660_ (.A(_1888_),
    .B(_1889_),
    .X(_1890_));
 sky130_fd_sc_hd__a21o_1 _5661_ (.A1(_1660_),
    .A2(_1865_),
    .B1(_1890_),
    .X(_1891_));
 sky130_fd_sc_hd__nand3_1 _5662_ (.A(_1660_),
    .B(_1865_),
    .C(_1890_),
    .Y(_1892_));
 sky130_fd_sc_hd__and2_1 _5663_ (.A(_1891_),
    .B(_1892_),
    .X(_1894_));
 sky130_fd_sc_hd__a31oi_2 _5664_ (.A1(_1029_),
    .A2(_0684_),
    .A3(_1668_),
    .B1(_1666_),
    .Y(_1895_));
 sky130_fd_sc_hd__xnor2_1 _5665_ (.A(_1894_),
    .B(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__o21a_1 _5666_ (.A1(_1863_),
    .A2(_1864_),
    .B1(_1896_),
    .X(_1897_));
 sky130_fd_sc_hd__or3_1 _5667_ (.A(_1863_),
    .B(_1864_),
    .C(_1896_),
    .X(_1898_));
 sky130_fd_sc_hd__and2b_1 _5668_ (.A_N(_1897_),
    .B(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__nor2_1 _5669_ (.A(_1681_),
    .B(_1684_),
    .Y(_1900_));
 sky130_fd_sc_hd__xnor2_2 _5670_ (.A(_1899_),
    .B(_1900_),
    .Y(_1901_));
 sky130_fd_sc_hd__and2_1 _5671_ (.A(_1790_),
    .B(_1801_),
    .X(_1902_));
 sky130_fd_sc_hd__and2b_1 _5672_ (.A_N(_1785_),
    .B(_1787_),
    .X(_1903_));
 sky130_fd_sc_hd__and2b_1 _5673_ (.A_N(_1788_),
    .B(_1749_),
    .X(_1905_));
 sky130_fd_sc_hd__nand2_1 _5674_ (.A(_1750_),
    .B(_1759_),
    .Y(_1906_));
 sky130_fd_sc_hd__nand2_1 _5675_ (.A(_1602_),
    .B(_2859_),
    .Y(_1907_));
 sky130_fd_sc_hd__nand2_1 _5676_ (.A(_1602_),
    .B(_2445_),
    .Y(_1908_));
 sky130_fd_sc_hd__and3_1 _5677_ (.A(_1229_),
    .B(_2858_),
    .C(_1908_),
    .X(_1909_));
 sky130_fd_sc_hd__xor2_1 _5678_ (.A(_1907_),
    .B(_1909_),
    .X(_1910_));
 sky130_fd_sc_hd__o21a_1 _5679_ (.A1(_0399_),
    .A2(_1758_),
    .B1(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__nor3_1 _5680_ (.A(_0399_),
    .B(_1758_),
    .C(_1910_),
    .Y(_1912_));
 sky130_fd_sc_hd__or2_1 _5681_ (.A(_1911_),
    .B(_1912_),
    .X(_1913_));
 sky130_fd_sc_hd__nand2_1 _5682_ (.A(_0388_),
    .B(_2845_),
    .Y(_1914_));
 sky130_fd_sc_hd__a21oi_1 _5683_ (.A1(_1752_),
    .A2(_1754_),
    .B1(_1757_),
    .Y(_1916_));
 sky130_fd_sc_hd__xnor2_1 _5684_ (.A(_1914_),
    .B(_1916_),
    .Y(_1917_));
 sky130_fd_sc_hd__nor2_1 _5685_ (.A(_1913_),
    .B(_1917_),
    .Y(_1918_));
 sky130_fd_sc_hd__and2_1 _5686_ (.A(_1913_),
    .B(_1917_),
    .X(_1919_));
 sky130_fd_sc_hd__or2_1 _5687_ (.A(_1918_),
    .B(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__a21o_1 _5688_ (.A1(_1906_),
    .A2(_1770_),
    .B1(_1920_),
    .X(_1921_));
 sky130_fd_sc_hd__nand3_1 _5689_ (.A(_1906_),
    .B(_1770_),
    .C(_1920_),
    .Y(_1922_));
 sky130_fd_sc_hd__nand2_1 _5690_ (.A(_1921_),
    .B(_1922_),
    .Y(_1923_));
 sky130_fd_sc_hd__nand2_1 _5691_ (.A(_0079_),
    .B(_2551_),
    .Y(_1924_));
 sky130_fd_sc_hd__o21ai_1 _5692_ (.A1(_1764_),
    .A2(_1767_),
    .B1(_1765_),
    .Y(_1925_));
 sky130_fd_sc_hd__xnor2_1 _5693_ (.A(_1924_),
    .B(_1925_),
    .Y(_1927_));
 sky130_fd_sc_hd__xnor2_1 _5694_ (.A(_1923_),
    .B(_1927_),
    .Y(_1928_));
 sky130_fd_sc_hd__a32o_1 _5695_ (.A1(_1770_),
    .A2(_1771_),
    .A3(_1775_),
    .B1(_1776_),
    .B2(_1783_),
    .X(_1929_));
 sky130_fd_sc_hd__xnor2_1 _5696_ (.A(_1928_),
    .B(_1929_),
    .Y(_1930_));
 sky130_fd_sc_hd__a31oi_2 _5697_ (.A1(_1029_),
    .A2(_2676_),
    .A3(_1781_),
    .B1(_1779_),
    .Y(_1931_));
 sky130_fd_sc_hd__xnor2_1 _5698_ (.A(_1930_),
    .B(_1931_),
    .Y(_1932_));
 sky130_fd_sc_hd__o21ai_1 _5699_ (.A1(_1903_),
    .A2(_1905_),
    .B1(_1932_),
    .Y(_1933_));
 sky130_fd_sc_hd__nor3_2 _5700_ (.A(_1903_),
    .B(_1905_),
    .C(_1932_),
    .Y(_1934_));
 sky130_fd_sc_hd__inv_2 _5701_ (.A(_1934_),
    .Y(_1935_));
 sky130_fd_sc_hd__nand2_1 _5702_ (.A(_1933_),
    .B(_1935_),
    .Y(_1936_));
 sky130_fd_sc_hd__or2_1 _5703_ (.A(_1902_),
    .B(_1936_),
    .X(_1938_));
 sky130_fd_sc_hd__nand2_1 _5704_ (.A(_1902_),
    .B(_1936_),
    .Y(_1939_));
 sky130_fd_sc_hd__and3_1 _5705_ (.A(_2885_),
    .B(_1938_),
    .C(_1939_),
    .X(_1940_));
 sky130_fd_sc_hd__and2b_1 _5706_ (.A_N(_1733_),
    .B(_1731_),
    .X(_1941_));
 sky130_fd_sc_hd__inv_2 _5707_ (.A(_1941_),
    .Y(_1942_));
 sky130_fd_sc_hd__or2b_1 _5708_ (.A(_1690_),
    .B_N(_1730_),
    .X(_1943_));
 sky130_fd_sc_hd__and3_1 _5709_ (.A(_1712_),
    .B(_1713_),
    .C(_1716_),
    .X(_1944_));
 sky130_fd_sc_hd__nor2_1 _5710_ (.A(_1717_),
    .B(_1725_),
    .Y(_1945_));
 sky130_fd_sc_hd__nand2_1 _5711_ (.A(_1693_),
    .B(_1702_),
    .Y(_1946_));
 sky130_fd_sc_hd__nand2_1 _5712_ (.A(_0698_),
    .B(_0530_),
    .Y(_1947_));
 sky130_fd_sc_hd__nand2_1 _5713_ (.A(_0573_),
    .B(_0530_),
    .Y(_1949_));
 sky130_fd_sc_hd__and3_1 _5714_ (.A(_0697_),
    .B(_2862_),
    .C(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__xor2_1 _5715_ (.A(_1947_),
    .B(_1950_),
    .X(_1951_));
 sky130_fd_sc_hd__xnor2_1 _5716_ (.A(_1700_),
    .B(_1951_),
    .Y(_1952_));
 sky130_fd_sc_hd__and3_1 _5717_ (.A(_2856_),
    .B(_0569_),
    .C(_1697_),
    .X(_1953_));
 sky130_fd_sc_hd__o21ba_1 _5718_ (.A1(_0704_),
    .A2(_1698_),
    .B1_N(_1953_),
    .X(_1954_));
 sky130_fd_sc_hd__xnor2_1 _5719_ (.A(_1708_),
    .B(_1954_),
    .Y(_1955_));
 sky130_fd_sc_hd__or2_1 _5720_ (.A(_1952_),
    .B(_1955_),
    .X(_1956_));
 sky130_fd_sc_hd__nand2_1 _5721_ (.A(_1952_),
    .B(_1955_),
    .Y(_1957_));
 sky130_fd_sc_hd__nand2_1 _5722_ (.A(_1956_),
    .B(_1957_),
    .Y(_1958_));
 sky130_fd_sc_hd__a21o_1 _5723_ (.A1(_1946_),
    .A2(_1712_),
    .B1(_1958_),
    .X(_1960_));
 sky130_fd_sc_hd__nand3_1 _5724_ (.A(_1946_),
    .B(_1712_),
    .C(_1958_),
    .Y(_1961_));
 sky130_fd_sc_hd__nand2_1 _5725_ (.A(_1960_),
    .B(_1961_),
    .Y(_1962_));
 sky130_fd_sc_hd__nor2_1 _5726_ (.A(_0545_),
    .B(_1708_),
    .Y(_1963_));
 sky130_fd_sc_hd__o21ai_1 _5727_ (.A1(_1706_),
    .A2(_1963_),
    .B1(_1709_),
    .Y(_1964_));
 sky130_fd_sc_hd__and3b_1 _5728_ (.A_N(_1964_),
    .B(_0674_),
    .C(_0546_),
    .X(_1965_));
 sky130_fd_sc_hd__a21bo_1 _5729_ (.A1(_0546_),
    .A2(_0685_),
    .B1_N(_1964_),
    .X(_1966_));
 sky130_fd_sc_hd__or2b_1 _5730_ (.A(_1965_),
    .B_N(_1966_),
    .X(_1967_));
 sky130_fd_sc_hd__xor2_1 _5731_ (.A(_1962_),
    .B(_1967_),
    .X(_1968_));
 sky130_fd_sc_hd__o21ai_1 _5732_ (.A1(_1944_),
    .A2(_1945_),
    .B1(_1968_),
    .Y(_1969_));
 sky130_fd_sc_hd__or3_1 _5733_ (.A(_1944_),
    .B(_1945_),
    .C(_1968_),
    .X(_1971_));
 sky130_fd_sc_hd__and2_1 _5734_ (.A(_1969_),
    .B(_1971_),
    .X(_1972_));
 sky130_fd_sc_hd__a31o_1 _5735_ (.A1(_0684_),
    .A2(_0696_),
    .A3(_1723_),
    .B1(_1721_),
    .X(_1973_));
 sky130_fd_sc_hd__xnor2_1 _5736_ (.A(_1972_),
    .B(_1973_),
    .Y(_1974_));
 sky130_fd_sc_hd__a21oi_2 _5737_ (.A1(_1727_),
    .A2(_1943_),
    .B1(_1974_),
    .Y(_1975_));
 sky130_fd_sc_hd__inv_2 _5738_ (.A(_1975_),
    .Y(_1976_));
 sky130_fd_sc_hd__nand3_2 _5739_ (.A(_1727_),
    .B(_1943_),
    .C(_1974_),
    .Y(_1977_));
 sky130_fd_sc_hd__nand2_1 _5740_ (.A(_1976_),
    .B(_1977_),
    .Y(_1978_));
 sky130_fd_sc_hd__a21oi_1 _5741_ (.A1(_1942_),
    .A2(_1742_),
    .B1(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__nand2_2 _5742_ (.A(_2882_),
    .B(_2883_),
    .Y(_1980_));
 sky130_fd_sc_hd__a31o_1 _5743_ (.A1(_1942_),
    .A2(_1742_),
    .A3(_1978_),
    .B1(_1980_),
    .X(_1982_));
 sky130_fd_sc_hd__nor2_1 _5744_ (.A(_1979_),
    .B(_1982_),
    .Y(_1983_));
 sky130_fd_sc_hd__clkinv_2 _5745_ (.A(_2878_),
    .Y(_1984_));
 sky130_fd_sc_hd__and2b_1 _5746_ (.A_N(_1841_),
    .B(_1843_),
    .X(_1985_));
 sky130_fd_sc_hd__and2b_1 _5747_ (.A_N(_1844_),
    .B(_1805_),
    .X(_1986_));
 sky130_fd_sc_hd__nand2_1 _5748_ (.A(_1807_),
    .B(_1815_),
    .Y(_1987_));
 sky130_fd_sc_hd__nand2_1 _5749_ (.A(_2859_),
    .B(_0530_),
    .Y(_1988_));
 sky130_fd_sc_hd__nand2_1 _5750_ (.A(_0530_),
    .B(_2445_),
    .Y(_1989_));
 sky130_fd_sc_hd__and3_1 _5751_ (.A(_2858_),
    .B(_2862_),
    .C(_1989_),
    .X(_1990_));
 sky130_fd_sc_hd__xor2_1 _5752_ (.A(_1988_),
    .B(_1990_),
    .X(_1991_));
 sky130_fd_sc_hd__o21a_1 _5753_ (.A1(_2857_),
    .A2(_1814_),
    .B1(_1991_),
    .X(_1993_));
 sky130_fd_sc_hd__nor3_1 _5754_ (.A(_2857_),
    .B(_1814_),
    .C(_1991_),
    .Y(_1994_));
 sky130_fd_sc_hd__or2_1 _5755_ (.A(_1993_),
    .B(_1994_),
    .X(_1995_));
 sky130_fd_sc_hd__nand2_1 _5756_ (.A(_2845_),
    .B(_2833_),
    .Y(_1996_));
 sky130_fd_sc_hd__a21oi_1 _5757_ (.A1(_1808_),
    .A2(_1810_),
    .B1(_1813_),
    .Y(_1997_));
 sky130_fd_sc_hd__xnor2_1 _5758_ (.A(_1996_),
    .B(_1997_),
    .Y(_1998_));
 sky130_fd_sc_hd__nor2_1 _5759_ (.A(_1995_),
    .B(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__and2_1 _5760_ (.A(_1995_),
    .B(_1998_),
    .X(_2000_));
 sky130_fd_sc_hd__or2_1 _5761_ (.A(_1999_),
    .B(_2000_),
    .X(_2001_));
 sky130_fd_sc_hd__a21o_1 _5762_ (.A1(_1987_),
    .A2(_1826_),
    .B1(_2001_),
    .X(_2002_));
 sky130_fd_sc_hd__nand3_1 _5763_ (.A(_1987_),
    .B(_1826_),
    .C(_2001_),
    .Y(_2004_));
 sky130_fd_sc_hd__nand2_1 _5764_ (.A(_2002_),
    .B(_2004_),
    .Y(_2005_));
 sky130_fd_sc_hd__o21ai_1 _5765_ (.A1(_1820_),
    .A2(_1823_),
    .B1(_1821_),
    .Y(_2006_));
 sky130_fd_sc_hd__and3b_1 _5766_ (.A_N(_2006_),
    .B(_0685_),
    .C(_2551_),
    .X(_2007_));
 sky130_fd_sc_hd__a21bo_1 _5767_ (.A1(_2551_),
    .A2(_0685_),
    .B1_N(_2006_),
    .X(_2008_));
 sky130_fd_sc_hd__or2b_1 _5768_ (.A(_2007_),
    .B_N(_2008_),
    .X(_2009_));
 sky130_fd_sc_hd__xnor2_1 _5769_ (.A(_2005_),
    .B(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__a32o_1 _5770_ (.A1(_1826_),
    .A2(_1827_),
    .A3(_1831_),
    .B1(_1832_),
    .B2(_1840_),
    .X(_2011_));
 sky130_fd_sc_hd__xnor2_1 _5771_ (.A(_2010_),
    .B(_2011_),
    .Y(_2012_));
 sky130_fd_sc_hd__a31oi_2 _5772_ (.A1(_2676_),
    .A2(_0696_),
    .A3(_1837_),
    .B1(_1835_),
    .Y(_2013_));
 sky130_fd_sc_hd__xnor2_1 _5773_ (.A(_2012_),
    .B(_2013_),
    .Y(_2015_));
 sky130_fd_sc_hd__o21ai_2 _5774_ (.A1(_1985_),
    .A2(_1986_),
    .B1(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__nor3_2 _5775_ (.A(_1985_),
    .B(_1986_),
    .C(_2015_),
    .Y(_2017_));
 sky130_fd_sc_hd__inv_2 _5776_ (.A(_2017_),
    .Y(_2018_));
 sky130_fd_sc_hd__nand2_1 _5777_ (.A(_2016_),
    .B(_2018_),
    .Y(_2019_));
 sky130_fd_sc_hd__a21oi_1 _5778_ (.A1(_1846_),
    .A2(_1856_),
    .B1(_2019_),
    .Y(_2020_));
 sky130_fd_sc_hd__and3_1 _5779_ (.A(_1846_),
    .B(_1856_),
    .C(_2019_),
    .X(_2021_));
 sky130_fd_sc_hd__o31a_1 _5780_ (.A1(_1984_),
    .A2(_2020_),
    .A3(_2021_),
    .B1(_1627_),
    .X(_2022_));
 sky130_fd_sc_hd__or3b_1 _5781_ (.A(_1940_),
    .B(_1983_),
    .C_N(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__o211a_2 _5782_ (.A1(_1631_),
    .A2(_1901_),
    .B1(_2023_),
    .C1(_1862_),
    .X(net20));
 sky130_fd_sc_hd__and2b_1 _5783_ (.A_N(_0698_),
    .B(_0573_),
    .X(_2025_));
 sky130_fd_sc_hd__a21o_1 _5784_ (.A1(_1602_),
    .A2(_0697_),
    .B1(_0698_),
    .X(_2026_));
 sky130_fd_sc_hd__o211a_1 _5785_ (.A1(_1638_),
    .A2(_2025_),
    .B1(_2026_),
    .C1(_1229_),
    .X(_2027_));
 sky130_fd_sc_hd__o21ai_1 _5786_ (.A1(_1872_),
    .A2(_1877_),
    .B1(_2027_),
    .Y(_2028_));
 sky130_fd_sc_hd__or3_1 _5787_ (.A(_1872_),
    .B(_1877_),
    .C(_2027_),
    .X(_2029_));
 sky130_fd_sc_hd__nand2_1 _5788_ (.A(_2028_),
    .B(_2029_),
    .Y(_2030_));
 sky130_fd_sc_hd__nor2_1 _5789_ (.A(_1874_),
    .B(_1875_),
    .Y(_2031_));
 sky130_fd_sc_hd__and2_1 _5790_ (.A(_1029_),
    .B(_2031_),
    .X(_2032_));
 sky130_fd_sc_hd__a21oi_1 _5791_ (.A1(_1585_),
    .A2(_1029_),
    .B1(_2031_),
    .Y(_2033_));
 sky130_fd_sc_hd__nor2_1 _5792_ (.A(_2032_),
    .B(_2033_),
    .Y(_2034_));
 sky130_fd_sc_hd__xnor2_1 _5793_ (.A(_2030_),
    .B(_2034_),
    .Y(_2036_));
 sky130_fd_sc_hd__nor2_1 _5794_ (.A(_1880_),
    .B(_1888_),
    .Y(_2037_));
 sky130_fd_sc_hd__xnor2_1 _5795_ (.A(_2036_),
    .B(_2037_),
    .Y(_2038_));
 sky130_fd_sc_hd__nand2_1 _5796_ (.A(_1885_),
    .B(_2038_),
    .Y(_2039_));
 sky130_fd_sc_hd__or2_1 _5797_ (.A(_1885_),
    .B(_2038_),
    .X(_2040_));
 sky130_fd_sc_hd__nand2_1 _5798_ (.A(_2039_),
    .B(_2040_),
    .Y(_2041_));
 sky130_fd_sc_hd__or2b_1 _5799_ (.A(_1895_),
    .B_N(_1894_),
    .X(_2042_));
 sky130_fd_sc_hd__nand2_1 _5800_ (.A(_1891_),
    .B(_2042_),
    .Y(_2043_));
 sky130_fd_sc_hd__xnor2_2 _5801_ (.A(_2041_),
    .B(_2043_),
    .Y(_2044_));
 sky130_fd_sc_hd__o31a_1 _5802_ (.A1(_1681_),
    .A2(_1684_),
    .A3(_1897_),
    .B1(_1898_),
    .X(_2045_));
 sky130_fd_sc_hd__xor2_2 _5803_ (.A(_2044_),
    .B(_2045_),
    .X(_2047_));
 sky130_fd_sc_hd__and2_1 _5804_ (.A(_1790_),
    .B(_1933_),
    .X(_2048_));
 sky130_fd_sc_hd__nor2_1 _5805_ (.A(_1924_),
    .B(_1925_),
    .Y(_2049_));
 sky130_fd_sc_hd__and2b_1 _5806_ (.A_N(_2859_),
    .B(_2445_),
    .X(_2050_));
 sky130_fd_sc_hd__a21o_1 _5807_ (.A1(_1602_),
    .A2(_2858_),
    .B1(_2859_),
    .X(_2051_));
 sky130_fd_sc_hd__o211a_1 _5808_ (.A1(_1753_),
    .A2(_2050_),
    .B1(_2051_),
    .C1(_1229_),
    .X(_2052_));
 sky130_fd_sc_hd__o21ai_1 _5809_ (.A1(_1912_),
    .A2(_1918_),
    .B1(_2052_),
    .Y(_2053_));
 sky130_fd_sc_hd__or3_1 _5810_ (.A(_1912_),
    .B(_1918_),
    .C(_2052_),
    .X(_2054_));
 sky130_fd_sc_hd__nand2_1 _5811_ (.A(_2053_),
    .B(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__nor2_1 _5812_ (.A(_1914_),
    .B(_1916_),
    .Y(_2056_));
 sky130_fd_sc_hd__and2_1 _5813_ (.A(_0079_),
    .B(_2056_),
    .X(_2058_));
 sky130_fd_sc_hd__a21oi_1 _5814_ (.A1(_0079_),
    .A2(_2845_),
    .B1(_2056_),
    .Y(_2059_));
 sky130_fd_sc_hd__nor2_1 _5815_ (.A(_2058_),
    .B(_2059_),
    .Y(_2060_));
 sky130_fd_sc_hd__xnor2_1 _5816_ (.A(_2055_),
    .B(_2060_),
    .Y(_2061_));
 sky130_fd_sc_hd__o21a_1 _5817_ (.A1(_1923_),
    .A2(_1927_),
    .B1(_1921_),
    .X(_2062_));
 sky130_fd_sc_hd__xnor2_1 _5818_ (.A(_2061_),
    .B(_2062_),
    .Y(_2063_));
 sky130_fd_sc_hd__nand2_1 _5819_ (.A(_2049_),
    .B(_2063_),
    .Y(_2064_));
 sky130_fd_sc_hd__or2_1 _5820_ (.A(_2049_),
    .B(_2063_),
    .X(_2065_));
 sky130_fd_sc_hd__nand2_1 _5821_ (.A(_2064_),
    .B(_2065_),
    .Y(_2066_));
 sky130_fd_sc_hd__or2b_1 _5822_ (.A(_1928_),
    .B_N(_1929_),
    .X(_2067_));
 sky130_fd_sc_hd__or2b_1 _5823_ (.A(_1931_),
    .B_N(_1930_),
    .X(_2069_));
 sky130_fd_sc_hd__nand2_1 _5824_ (.A(_2067_),
    .B(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__xor2_1 _5825_ (.A(_2066_),
    .B(_2070_),
    .X(_2071_));
 sky130_fd_sc_hd__a211o_1 _5826_ (.A1(_1801_),
    .A2(_2048_),
    .B1(_2071_),
    .C1(_1934_),
    .X(_2072_));
 sky130_fd_sc_hd__a21o_1 _5827_ (.A1(_1801_),
    .A2(_2048_),
    .B1(_1934_),
    .X(_2073_));
 sky130_fd_sc_hd__nand2_1 _5828_ (.A(_2071_),
    .B(_2073_),
    .Y(_2074_));
 sky130_fd_sc_hd__a21o_1 _5829_ (.A1(_2858_),
    .A2(_0530_),
    .B1(_2859_),
    .X(_2075_));
 sky130_fd_sc_hd__o211a_1 _5830_ (.A1(_1809_),
    .A2(_2050_),
    .B1(_2075_),
    .C1(_2862_),
    .X(_2076_));
 sky130_fd_sc_hd__o21ai_1 _5831_ (.A1(_1994_),
    .A2(_1999_),
    .B1(_2076_),
    .Y(_2077_));
 sky130_fd_sc_hd__or3_1 _5832_ (.A(_1994_),
    .B(_1999_),
    .C(_2076_),
    .X(_2078_));
 sky130_fd_sc_hd__nand2_1 _5833_ (.A(_2077_),
    .B(_2078_),
    .Y(_2080_));
 sky130_fd_sc_hd__nor2_1 _5834_ (.A(_1996_),
    .B(_1997_),
    .Y(_2081_));
 sky130_fd_sc_hd__and2_1 _5835_ (.A(_0685_),
    .B(_2081_),
    .X(_2082_));
 sky130_fd_sc_hd__a21oi_1 _5836_ (.A1(_2845_),
    .A2(_0696_),
    .B1(_2081_),
    .Y(_2083_));
 sky130_fd_sc_hd__nor2_1 _5837_ (.A(_2082_),
    .B(_2083_),
    .Y(_2084_));
 sky130_fd_sc_hd__xnor2_1 _5838_ (.A(_2080_),
    .B(_2084_),
    .Y(_2085_));
 sky130_fd_sc_hd__o21a_1 _5839_ (.A1(_2005_),
    .A2(_2009_),
    .B1(_2002_),
    .X(_2086_));
 sky130_fd_sc_hd__xnor2_1 _5840_ (.A(_2085_),
    .B(_2086_),
    .Y(_2087_));
 sky130_fd_sc_hd__nand2_1 _5841_ (.A(_2007_),
    .B(_2087_),
    .Y(_2088_));
 sky130_fd_sc_hd__or2_1 _5842_ (.A(_2007_),
    .B(_2087_),
    .X(_2089_));
 sky130_fd_sc_hd__nand2_1 _5843_ (.A(_2088_),
    .B(_2089_),
    .Y(_2091_));
 sky130_fd_sc_hd__or2b_1 _5844_ (.A(_2010_),
    .B_N(_2011_),
    .X(_2092_));
 sky130_fd_sc_hd__or2b_1 _5845_ (.A(_2013_),
    .B_N(_2012_),
    .X(_2093_));
 sky130_fd_sc_hd__nand2_1 _5846_ (.A(_2092_),
    .B(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hd__xor2_1 _5847_ (.A(_2091_),
    .B(_2094_),
    .X(_2095_));
 sky130_fd_sc_hd__a31o_1 _5848_ (.A1(_1846_),
    .A2(_1856_),
    .A3(_2016_),
    .B1(_2017_),
    .X(_2096_));
 sky130_fd_sc_hd__xor2_1 _5849_ (.A(_2095_),
    .B(_2096_),
    .X(_2097_));
 sky130_fd_sc_hd__a32o_1 _5850_ (.A1(_2885_),
    .A2(_2072_),
    .A3(_2074_),
    .B1(_2879_),
    .B2(_2097_),
    .X(_2098_));
 sky130_fd_sc_hd__nand2_1 _5851_ (.A(_1972_),
    .B(_1973_),
    .Y(_2099_));
 sky130_fd_sc_hd__o21ai_1 _5852_ (.A1(_1700_),
    .A2(_1951_),
    .B1(_1956_),
    .Y(_2100_));
 sky130_fd_sc_hd__a21o_1 _5853_ (.A1(_0697_),
    .A2(_0530_),
    .B1(_0698_),
    .X(_2102_));
 sky130_fd_sc_hd__o211a_1 _5854_ (.A1(_1695_),
    .A2(_2025_),
    .B1(_2102_),
    .C1(_2862_),
    .X(_2103_));
 sky130_fd_sc_hd__xnor2_1 _5855_ (.A(_2100_),
    .B(_2103_),
    .Y(_2104_));
 sky130_fd_sc_hd__nor2_1 _5856_ (.A(_1708_),
    .B(_1954_),
    .Y(_2105_));
 sky130_fd_sc_hd__and2_1 _5857_ (.A(_0685_),
    .B(_2105_),
    .X(_2106_));
 sky130_fd_sc_hd__a21oi_1 _5858_ (.A1(_1585_),
    .A2(_0696_),
    .B1(_2105_),
    .Y(_2107_));
 sky130_fd_sc_hd__nor2_1 _5859_ (.A(_2106_),
    .B(_2107_),
    .Y(_2108_));
 sky130_fd_sc_hd__xnor2_1 _5860_ (.A(_2104_),
    .B(_2108_),
    .Y(_2109_));
 sky130_fd_sc_hd__o21a_1 _5861_ (.A1(_1962_),
    .A2(_1967_),
    .B1(_1960_),
    .X(_2110_));
 sky130_fd_sc_hd__xnor2_1 _5862_ (.A(_2109_),
    .B(_2110_),
    .Y(_2111_));
 sky130_fd_sc_hd__nand2_1 _5863_ (.A(_1965_),
    .B(_2111_),
    .Y(_2113_));
 sky130_fd_sc_hd__or2_1 _5864_ (.A(_1965_),
    .B(_2111_),
    .X(_2114_));
 sky130_fd_sc_hd__nand2_1 _5865_ (.A(_2113_),
    .B(_2114_),
    .Y(_2115_));
 sky130_fd_sc_hd__a21o_1 _5866_ (.A1(_1969_),
    .A2(_2099_),
    .B1(_2115_),
    .X(_2116_));
 sky130_fd_sc_hd__nand3_1 _5867_ (.A(_1969_),
    .B(_2099_),
    .C(_2115_),
    .Y(_2117_));
 sky130_fd_sc_hd__nand2_1 _5868_ (.A(_2116_),
    .B(_2117_),
    .Y(_2118_));
 sky130_fd_sc_hd__inv_2 _5869_ (.A(_1977_),
    .Y(_2119_));
 sky130_fd_sc_hd__a31o_1 _5870_ (.A1(_1942_),
    .A2(_1742_),
    .A3(_1976_),
    .B1(_2119_),
    .X(_2120_));
 sky130_fd_sc_hd__a311o_1 _5871_ (.A1(_1942_),
    .A2(_1742_),
    .A3(_1976_),
    .B1(_2119_),
    .C1(_2118_),
    .X(_2121_));
 sky130_fd_sc_hd__nand2_1 _5872_ (.A(_1744_),
    .B(_2121_),
    .Y(_2122_));
 sky130_fd_sc_hd__a21o_1 _5873_ (.A1(_2118_),
    .A2(_2120_),
    .B1(_2122_),
    .X(_2124_));
 sky130_fd_sc_hd__or3b_1 _5874_ (.A(_1025_),
    .B(_2098_),
    .C_N(_2124_),
    .X(_2125_));
 sky130_fd_sc_hd__o211a_2 _5875_ (.A1(_1631_),
    .A2(_2047_),
    .B1(_2125_),
    .C1(_1862_),
    .X(net21));
 sky130_fd_sc_hd__and3_1 _5876_ (.A(_2039_),
    .B(_2040_),
    .C(_2043_),
    .X(_2126_));
 sky130_fd_sc_hd__o311a_1 _5877_ (.A1(_1681_),
    .A2(_1684_),
    .A3(_1897_),
    .B1(_1898_),
    .C1(_2044_),
    .X(_2127_));
 sky130_fd_sc_hd__o21ai_1 _5878_ (.A1(_1880_),
    .A2(_1888_),
    .B1(_2036_),
    .Y(_2128_));
 sky130_fd_sc_hd__or2b_1 _5879_ (.A(_2030_),
    .B_N(_2034_),
    .X(_2129_));
 sky130_fd_sc_hd__nand4_1 _5880_ (.A(_0698_),
    .B(_1602_),
    .C(_0697_),
    .D(_1229_),
    .Y(_2130_));
 sky130_fd_sc_hd__a21oi_1 _5881_ (.A1(_2028_),
    .A2(_2129_),
    .B1(_2130_),
    .Y(_2131_));
 sky130_fd_sc_hd__and3_1 _5882_ (.A(_2028_),
    .B(_2129_),
    .C(_2130_),
    .X(_2132_));
 sky130_fd_sc_hd__nor2_1 _5883_ (.A(_2131_),
    .B(_2132_),
    .Y(_2134_));
 sky130_fd_sc_hd__xnor2_1 _5884_ (.A(_2032_),
    .B(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__a21oi_1 _5885_ (.A1(_2128_),
    .A2(_2039_),
    .B1(_2135_),
    .Y(_2136_));
 sky130_fd_sc_hd__and3_1 _5886_ (.A(_2128_),
    .B(_2039_),
    .C(_2135_),
    .X(_2137_));
 sky130_fd_sc_hd__nor2_1 _5887_ (.A(_2136_),
    .B(_2137_),
    .Y(_2138_));
 sky130_fd_sc_hd__nor3b_2 _5888_ (.A(_2126_),
    .B(_2127_),
    .C_N(_2138_),
    .Y(_2139_));
 sky130_fd_sc_hd__o21ba_1 _5889_ (.A1(_2126_),
    .A2(_2127_),
    .B1_N(_2138_),
    .X(_2140_));
 sky130_fd_sc_hd__or2b_1 _5890_ (.A(_2091_),
    .B_N(_2094_),
    .X(_2141_));
 sky130_fd_sc_hd__a311o_1 _5891_ (.A1(_1846_),
    .A2(_1856_),
    .A3(_2016_),
    .B1(_2017_),
    .C1(_2095_),
    .X(_2142_));
 sky130_fd_sc_hd__or2b_1 _5892_ (.A(_2086_),
    .B_N(_2085_),
    .X(_2143_));
 sky130_fd_sc_hd__nand4_2 _5893_ (.A(_2859_),
    .B(_2858_),
    .C(_0530_),
    .D(_2862_),
    .Y(_2145_));
 sky130_fd_sc_hd__or2b_1 _5894_ (.A(_2080_),
    .B_N(_2084_),
    .X(_2146_));
 sky130_fd_sc_hd__nand2_1 _5895_ (.A(_2077_),
    .B(_2146_),
    .Y(_2147_));
 sky130_fd_sc_hd__xnor2_1 _5896_ (.A(_2145_),
    .B(_2147_),
    .Y(_2148_));
 sky130_fd_sc_hd__xnor2_1 _5897_ (.A(_2082_),
    .B(_2148_),
    .Y(_2149_));
 sky130_fd_sc_hd__a21oi_1 _5898_ (.A1(_2143_),
    .A2(_2088_),
    .B1(_2149_),
    .Y(_2150_));
 sky130_fd_sc_hd__and3_1 _5899_ (.A(_2143_),
    .B(_2088_),
    .C(_2149_),
    .X(_2151_));
 sky130_fd_sc_hd__or2_1 _5900_ (.A(_2150_),
    .B(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__nand3_1 _5901_ (.A(_2141_),
    .B(_2142_),
    .C(_2152_),
    .Y(_2153_));
 sky130_fd_sc_hd__a21o_1 _5902_ (.A1(_2141_),
    .A2(_2142_),
    .B1(_2152_),
    .X(_2154_));
 sky130_fd_sc_hd__and3_1 _5903_ (.A(_2879_),
    .B(_2153_),
    .C(_2154_),
    .X(_2156_));
 sky130_fd_sc_hd__or2b_1 _5904_ (.A(_2066_),
    .B_N(_2070_),
    .X(_2157_));
 sky130_fd_sc_hd__or2b_1 _5905_ (.A(_2062_),
    .B_N(_2061_),
    .X(_2158_));
 sky130_fd_sc_hd__nand4_1 _5906_ (.A(_1602_),
    .B(_1229_),
    .C(_2859_),
    .D(_2858_),
    .Y(_2159_));
 sky130_fd_sc_hd__or2b_1 _5907_ (.A(_2055_),
    .B_N(_2060_),
    .X(_2160_));
 sky130_fd_sc_hd__nand2_1 _5908_ (.A(_2053_),
    .B(_2160_),
    .Y(_2161_));
 sky130_fd_sc_hd__xnor2_1 _5909_ (.A(_2159_),
    .B(_2161_),
    .Y(_2162_));
 sky130_fd_sc_hd__xnor2_1 _5910_ (.A(_2058_),
    .B(_2162_),
    .Y(_2163_));
 sky130_fd_sc_hd__a21oi_2 _5911_ (.A1(_2158_),
    .A2(_2064_),
    .B1(_2163_),
    .Y(_2164_));
 sky130_fd_sc_hd__and3_1 _5912_ (.A(_2158_),
    .B(_2064_),
    .C(_2163_),
    .X(_2165_));
 sky130_fd_sc_hd__nor2_1 _5913_ (.A(_2164_),
    .B(_2165_),
    .Y(_2167_));
 sky130_fd_sc_hd__inv_2 _5914_ (.A(_2167_),
    .Y(_2168_));
 sky130_fd_sc_hd__nand3_1 _5915_ (.A(_2157_),
    .B(_2072_),
    .C(_2168_),
    .Y(_2169_));
 sky130_fd_sc_hd__a21o_1 _5916_ (.A1(_2157_),
    .A2(_2072_),
    .B1(_2168_),
    .X(_2170_));
 sky130_fd_sc_hd__and3_1 _5917_ (.A(_2884_),
    .B(_2169_),
    .C(_2170_),
    .X(_2171_));
 sky130_fd_sc_hd__or2b_1 _5918_ (.A(_2110_),
    .B_N(_2109_),
    .X(_2172_));
 sky130_fd_sc_hd__and4_1 _5919_ (.A(_0698_),
    .B(_0697_),
    .C(_0530_),
    .D(_2862_),
    .X(_2173_));
 sky130_fd_sc_hd__or2b_1 _5920_ (.A(_2104_),
    .B_N(_2108_),
    .X(_2174_));
 sky130_fd_sc_hd__a21bo_1 _5921_ (.A1(_2100_),
    .A2(_2103_),
    .B1_N(_2174_),
    .X(_2175_));
 sky130_fd_sc_hd__xor2_1 _5922_ (.A(_2173_),
    .B(_2175_),
    .X(_2176_));
 sky130_fd_sc_hd__or2_1 _5923_ (.A(_2106_),
    .B(_2176_),
    .X(_2178_));
 sky130_fd_sc_hd__nand2_1 _5924_ (.A(_2106_),
    .B(_2176_),
    .Y(_2179_));
 sky130_fd_sc_hd__nand2_1 _5925_ (.A(_2178_),
    .B(_2179_),
    .Y(_2180_));
 sky130_fd_sc_hd__a21oi_2 _5926_ (.A1(_2172_),
    .A2(_2113_),
    .B1(_2180_),
    .Y(_2181_));
 sky130_fd_sc_hd__and3_1 _5927_ (.A(_2172_),
    .B(_2113_),
    .C(_2180_),
    .X(_2182_));
 sky130_fd_sc_hd__or2_1 _5928_ (.A(_2181_),
    .B(_2182_),
    .X(_2183_));
 sky130_fd_sc_hd__a21oi_1 _5929_ (.A1(_2116_),
    .A2(_2121_),
    .B1(_2183_),
    .Y(_2184_));
 sky130_fd_sc_hd__a31o_1 _5930_ (.A1(_2116_),
    .A2(_2121_),
    .A3(_2183_),
    .B1(_1980_),
    .X(_2185_));
 sky130_fd_sc_hd__nor2_1 _5931_ (.A(_2184_),
    .B(_2185_),
    .Y(_2186_));
 sky130_fd_sc_hd__or4_1 _5932_ (.A(_1024_),
    .B(_2156_),
    .C(_2171_),
    .D(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__o311a_2 _5933_ (.A1(_1631_),
    .A2(_2139_),
    .A3(_2140_),
    .B1(_2187_),
    .C1(_1028_),
    .X(net22));
 sky130_fd_sc_hd__a211o_1 _5934_ (.A1(_2032_),
    .A2(_2134_),
    .B1(_2131_),
    .C1(_1627_),
    .X(_2189_));
 sky130_fd_sc_hd__inv_2 _5935_ (.A(_2137_),
    .Y(_2190_));
 sky130_fd_sc_hd__o31a_1 _5936_ (.A1(_2126_),
    .A2(_2127_),
    .A3(_2136_),
    .B1(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__a21oi_1 _5937_ (.A1(_2053_),
    .A2(_2160_),
    .B1(_2159_),
    .Y(_2192_));
 sky130_fd_sc_hd__a21oi_1 _5938_ (.A1(_2058_),
    .A2(_2162_),
    .B1(_2192_),
    .Y(_2193_));
 sky130_fd_sc_hd__inv_2 _5939_ (.A(_2164_),
    .Y(_2194_));
 sky130_fd_sc_hd__a31o_1 _5940_ (.A1(_2157_),
    .A2(_2072_),
    .A3(_2194_),
    .B1(_2165_),
    .X(_2195_));
 sky130_fd_sc_hd__a21bo_1 _5941_ (.A1(_2193_),
    .A2(_2195_),
    .B1_N(_2885_),
    .X(_2196_));
 sky130_fd_sc_hd__nand2_1 _5942_ (.A(_2173_),
    .B(_2175_),
    .Y(_2197_));
 sky130_fd_sc_hd__inv_2 _5943_ (.A(_2181_),
    .Y(_2199_));
 sky130_fd_sc_hd__a31o_1 _5944_ (.A1(_2116_),
    .A2(_2121_),
    .A3(_2199_),
    .B1(_2182_),
    .X(_2200_));
 sky130_fd_sc_hd__a41o_1 _5945_ (.A1(_2883_),
    .A2(_2197_),
    .A3(_2179_),
    .A4(_2200_),
    .B1(net15),
    .X(_2201_));
 sky130_fd_sc_hd__a21oi_1 _5946_ (.A1(_2077_),
    .A2(_2146_),
    .B1(_2145_),
    .Y(_2202_));
 sky130_fd_sc_hd__a21oi_1 _5947_ (.A1(_2082_),
    .A2(_2148_),
    .B1(_2202_),
    .Y(_2203_));
 sky130_fd_sc_hd__inv_2 _5948_ (.A(_2150_),
    .Y(_2204_));
 sky130_fd_sc_hd__a31o_1 _5949_ (.A1(_2141_),
    .A2(_2142_),
    .A3(_2204_),
    .B1(_2151_),
    .X(_2205_));
 sky130_fd_sc_hd__a21o_1 _5950_ (.A1(_2203_),
    .A2(_2205_),
    .B1(_1984_),
    .X(_2206_));
 sky130_fd_sc_hd__nand3_1 _5951_ (.A(_2196_),
    .B(_2201_),
    .C(_2206_),
    .Y(_2207_));
 sky130_fd_sc_hd__o211a_2 _5952_ (.A1(_2189_),
    .A2(_2191_),
    .B1(_2207_),
    .C1(_1862_),
    .X(net23));
 sky130_fd_sc_hd__a22o_1 _5953_ (.A1(_0964_),
    .A2(_2471_),
    .B1(_2778_),
    .B2(_0899_),
    .X(_2209_));
 sky130_fd_sc_hd__and3b_1 _5954_ (.A_N(_0978_),
    .B(_1744_),
    .C(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__a22o_1 _5955_ (.A1(_0280_),
    .A2(_2550_),
    .B1(_2717_),
    .B2(_0342_),
    .X(_2211_));
 sky130_fd_sc_hd__and3b_1 _5956_ (.A_N(_0345_),
    .B(_2885_),
    .C(_2211_),
    .X(_2212_));
 sky130_fd_sc_hd__inv_2 _5957_ (.A(_2796_),
    .Y(_2213_));
 sky130_fd_sc_hd__a22o_1 _5958_ (.A1(_2471_),
    .A2(_2550_),
    .B1(_2717_),
    .B2(_2778_),
    .X(_2214_));
 sky130_fd_sc_hd__a31o_1 _5959_ (.A1(_2213_),
    .A2(_2879_),
    .A3(_2214_),
    .B1(_1025_),
    .X(_2215_));
 sky130_fd_sc_hd__a22oi_1 _5960_ (.A1(_0280_),
    .A2(_0964_),
    .B1(_0342_),
    .B2(_0899_),
    .Y(_2216_));
 sky130_fd_sc_hd__o21ai_1 _5961_ (.A1(_1539_),
    .A2(_2216_),
    .B1(_1025_),
    .Y(_2217_));
 sky130_fd_sc_hd__o311a_1 _5962_ (.A1(_2210_),
    .A2(_2212_),
    .A3(_2215_),
    .B1(_2217_),
    .C1(_1028_),
    .X(net16));
 sky130_fd_sc_hd__and2_1 _5963_ (.A(_1540_),
    .B(_1541_),
    .X(_2219_));
 sky130_fd_sc_hd__nor2_1 _5964_ (.A(_1542_),
    .B(_2219_),
    .Y(_2220_));
 sky130_fd_sc_hd__and2_1 _5965_ (.A(_0979_),
    .B(_0980_),
    .X(_2221_));
 sky130_fd_sc_hd__nor2_1 _5966_ (.A(_0981_),
    .B(_2221_),
    .Y(_2222_));
 sky130_fd_sc_hd__a21bo_1 _5967_ (.A1(_0346_),
    .A2(_0347_),
    .B1_N(_2884_),
    .X(_2223_));
 sky130_fd_sc_hd__a21o_1 _5968_ (.A1(_2797_),
    .A2(_2798_),
    .B1(_1984_),
    .X(_2224_));
 sky130_fd_sc_hd__o22ai_1 _5969_ (.A1(_0348_),
    .A2(_2223_),
    .B1(_2224_),
    .B2(_2799_),
    .Y(_2225_));
 sky130_fd_sc_hd__a211o_1 _5970_ (.A1(_1744_),
    .A2(_2222_),
    .B1(_2225_),
    .C1(_1025_),
    .X(_2226_));
 sky130_fd_sc_hd__o211a_1 _5971_ (.A1(_1631_),
    .A2(_2220_),
    .B1(_2226_),
    .C1(_1862_),
    .X(net24));
 sky130_fd_sc_hd__and2_1 _5972_ (.A(_1536_),
    .B(_1544_),
    .X(_2227_));
 sky130_fd_sc_hd__nor2_1 _5973_ (.A(_1545_),
    .B(_2227_),
    .Y(_2229_));
 sky130_fd_sc_hd__o21ai_1 _5974_ (.A1(_2793_),
    .A2(_2800_),
    .B1(_2879_),
    .Y(_2230_));
 sky130_fd_sc_hd__o21a_1 _5975_ (.A1(_0341_),
    .A2(_0349_),
    .B1(_2884_),
    .X(_2231_));
 sky130_fd_sc_hd__and2_1 _5976_ (.A(_0972_),
    .B(_0975_),
    .X(_2232_));
 sky130_fd_sc_hd__o21ai_1 _5977_ (.A1(_2232_),
    .A2(_0983_),
    .B1(_1744_),
    .Y(_2233_));
 sky130_fd_sc_hd__o2bb2a_1 _5978_ (.A1_N(_2231_),
    .A2_N(_0350_),
    .B1(_0984_),
    .B2(_2233_),
    .X(_2234_));
 sky130_fd_sc_hd__o211ai_1 _5979_ (.A1(_2801_),
    .A2(_2230_),
    .B1(_2234_),
    .C1(_1631_),
    .Y(_2235_));
 sky130_fd_sc_hd__o211a_1 _5980_ (.A1(_1631_),
    .A2(_2229_),
    .B1(_2235_),
    .C1(_1862_),
    .X(net25));
 sky130_fd_sc_hd__o21ba_1 _5981_ (.A1(_1533_),
    .A2(_1534_),
    .B1_N(_1545_),
    .X(_2236_));
 sky130_fd_sc_hd__nor2_1 _5982_ (.A(_1546_),
    .B(_2236_),
    .Y(_2237_));
 sky130_fd_sc_hd__nand2_1 _5983_ (.A(_2791_),
    .B(_2801_),
    .Y(_2239_));
 sky130_fd_sc_hd__o21a_1 _5984_ (.A1(_2791_),
    .A2(_2801_),
    .B1(_2879_),
    .X(_2240_));
 sky130_fd_sc_hd__nand2_1 _5985_ (.A(_0974_),
    .B(_0984_),
    .Y(_2241_));
 sky130_fd_sc_hd__o21a_1 _5986_ (.A1(_0974_),
    .A2(_0984_),
    .B1(_1744_),
    .X(_2242_));
 sky130_fd_sc_hd__o21a_1 _5987_ (.A1(_0334_),
    .A2(_0339_),
    .B1(_0350_),
    .X(_2243_));
 sky130_fd_sc_hd__nor2_1 _5988_ (.A(_0351_),
    .B(_2243_),
    .Y(_2244_));
 sky130_fd_sc_hd__a22o_1 _5989_ (.A1(_2241_),
    .A2(_2242_),
    .B1(_2244_),
    .B2(_2885_),
    .X(_2245_));
 sky130_fd_sc_hd__a211o_1 _5990_ (.A1(_2239_),
    .A2(_2240_),
    .B1(_2245_),
    .C1(_1025_),
    .X(_2246_));
 sky130_fd_sc_hd__o211a_1 _5991_ (.A1(_1631_),
    .A2(_2237_),
    .B1(_2246_),
    .C1(_1862_),
    .X(net26));
 sky130_fd_sc_hd__xor2_1 _5992_ (.A(_0958_),
    .B(_0991_),
    .X(_2247_));
 sky130_fd_sc_hd__a21oi_1 _5993_ (.A1(_2241_),
    .A2(_2247_),
    .B1(_1980_),
    .Y(_2249_));
 sky130_fd_sc_hd__nor2_1 _5994_ (.A(_0338_),
    .B(_0334_),
    .Y(_2250_));
 sky130_fd_sc_hd__o21ba_1 _5995_ (.A1(_0335_),
    .A2(_2250_),
    .B1_N(_0351_),
    .X(_2251_));
 sky130_fd_sc_hd__or3_1 _5996_ (.A(_2882_),
    .B(_2883_),
    .C(_2251_),
    .X(_2252_));
 sky130_fd_sc_hd__a21oi_1 _5997_ (.A1(_2777_),
    .A2(_2787_),
    .B1(_2790_),
    .Y(_2253_));
 sky130_fd_sc_hd__or2_1 _5998_ (.A(_2788_),
    .B(_2253_),
    .X(_2254_));
 sky130_fd_sc_hd__a211o_1 _5999_ (.A1(_2239_),
    .A2(_2254_),
    .B1(_1984_),
    .C1(_2802_),
    .X(_2255_));
 sky130_fd_sc_hd__o211a_1 _6000_ (.A1(_0352_),
    .A2(_2252_),
    .B1(_2255_),
    .C1(_1627_),
    .X(_2256_));
 sky130_fd_sc_hd__a21bo_1 _6001_ (.A1(_0985_),
    .A2(_2249_),
    .B1_N(_2256_),
    .X(_2257_));
 sky130_fd_sc_hd__nor2_1 _6002_ (.A(_1533_),
    .B(_1546_),
    .Y(_2258_));
 sky130_fd_sc_hd__o21ai_1 _6003_ (.A1(_1518_),
    .A2(_2258_),
    .B1(_1024_),
    .Y(_2260_));
 sky130_fd_sc_hd__a21o_1 _6004_ (.A1(_1518_),
    .A2(_2258_),
    .B1(_2260_),
    .X(_2261_));
 sky130_fd_sc_hd__and3_1 _6005_ (.A(_1028_),
    .B(_2257_),
    .C(_2261_),
    .X(_2262_));
 sky130_fd_sc_hd__clkbuf_1 _6006_ (.A(_2262_),
    .X(net27));
 sky130_fd_sc_hd__or2_1 _6007_ (.A(_1550_),
    .B(_1551_),
    .X(_2263_));
 sky130_fd_sc_hd__xor2_1 _6008_ (.A(_1547_),
    .B(_2263_),
    .X(_2264_));
 sky130_fd_sc_hd__a21oi_1 _6009_ (.A1(_2803_),
    .A2(_2804_),
    .B1(_2802_),
    .Y(_2265_));
 sky130_fd_sc_hd__o21ai_1 _6010_ (.A1(_0988_),
    .A2(_0989_),
    .B1(_0985_),
    .Y(_2266_));
 sky130_fd_sc_hd__nand2_1 _6011_ (.A(_0352_),
    .B(_0354_),
    .Y(_2267_));
 sky130_fd_sc_hd__or2_1 _6012_ (.A(_0352_),
    .B(_0354_),
    .X(_2268_));
 sky130_fd_sc_hd__a31o_1 _6013_ (.A1(_2267_),
    .A2(_2885_),
    .A3(_2268_),
    .B1(_1024_),
    .X(_2270_));
 sky130_fd_sc_hd__a31oi_1 _6014_ (.A1(_0990_),
    .A2(_1744_),
    .A3(_2266_),
    .B1(_2270_),
    .Y(_2271_));
 sky130_fd_sc_hd__o31ai_1 _6015_ (.A1(_2805_),
    .A2(_1984_),
    .A3(_2265_),
    .B1(_2271_),
    .Y(_2272_));
 sky130_fd_sc_hd__o211a_1 _6016_ (.A1(_1631_),
    .A2(_2264_),
    .B1(_2272_),
    .C1(_1862_),
    .X(net28));
 sky130_fd_sc_hd__a211oi_1 _6017_ (.A1(_2773_),
    .A2(_2806_),
    .B1(_2789_),
    .C1(_2805_),
    .Y(_2273_));
 sky130_fd_sc_hd__and4b_1 _6018_ (.A_N(_2273_),
    .B(_2883_),
    .C(net15),
    .D(_2807_),
    .X(_2274_));
 sky130_fd_sc_hd__nor2_1 _6019_ (.A(_0355_),
    .B(_0359_),
    .Y(_2275_));
 sky130_fd_sc_hd__nand2_1 _6020_ (.A(_0355_),
    .B(_0359_),
    .Y(_2276_));
 sky130_fd_sc_hd__and3b_1 _6021_ (.A_N(_2275_),
    .B(_2884_),
    .C(_2276_),
    .X(_2277_));
 sky130_fd_sc_hd__nand2_1 _6022_ (.A(_0990_),
    .B(_0994_),
    .Y(_2278_));
 sky130_fd_sc_hd__nor2_1 _6023_ (.A(_0996_),
    .B(_0997_),
    .Y(_2280_));
 sky130_fd_sc_hd__xnor2_1 _6024_ (.A(_2278_),
    .B(_2280_),
    .Y(_2281_));
 sky130_fd_sc_hd__nor2_1 _6025_ (.A(_1980_),
    .B(_2281_),
    .Y(_2282_));
 sky130_fd_sc_hd__or3_1 _6026_ (.A(_1024_),
    .B(_2277_),
    .C(_2282_),
    .X(_2283_));
 sky130_fd_sc_hd__and2b_1 _6027_ (.A_N(_1559_),
    .B(_1558_),
    .X(_2284_));
 sky130_fd_sc_hd__xnor2_1 _6028_ (.A(_1555_),
    .B(_2284_),
    .Y(_2285_));
 sky130_fd_sc_hd__nand2_1 _6029_ (.A(_1025_),
    .B(_2285_),
    .Y(_2286_));
 sky130_fd_sc_hd__o211a_1 _6030_ (.A1(_2274_),
    .A2(_2283_),
    .B1(_2286_),
    .C1(_1862_),
    .X(net29));
 sky130_fd_sc_hd__and3_1 _6031_ (.A(_0270_),
    .B(_0271_),
    .C(_0307_),
    .X(_2287_));
 sky130_fd_sc_hd__nor2_1 _6032_ (.A(_0308_),
    .B(_2287_),
    .Y(_2288_));
 sky130_fd_sc_hd__o21ai_1 _6033_ (.A1(_0357_),
    .A2(_2275_),
    .B1(_2288_),
    .Y(_2290_));
 sky130_fd_sc_hd__or3_1 _6034_ (.A(_0357_),
    .B(_2275_),
    .C(_2288_),
    .X(_2291_));
 sky130_fd_sc_hd__and3b_1 _6035_ (.A_N(_2883_),
    .B(_2290_),
    .C(_2291_),
    .X(_2292_));
 sky130_fd_sc_hd__and3_1 _6036_ (.A(_2808_),
    .B(_2809_),
    .C(_2756_),
    .X(_2293_));
 sky130_fd_sc_hd__nor2_1 _6037_ (.A(_2810_),
    .B(_2293_),
    .Y(_2294_));
 sky130_fd_sc_hd__and2_1 _6038_ (.A(_2773_),
    .B(_2807_),
    .X(_2295_));
 sky130_fd_sc_hd__xnor2_1 _6039_ (.A(_2294_),
    .B(_2295_),
    .Y(_2296_));
 sky130_fd_sc_hd__and3_1 _6040_ (.A(_0908_),
    .B(_0909_),
    .C(_0943_),
    .X(_2297_));
 sky130_fd_sc_hd__nor2_1 _6041_ (.A(_0944_),
    .B(_2297_),
    .Y(_2298_));
 sky130_fd_sc_hd__and2b_1 _6042_ (.A_N(_0996_),
    .B(_0998_),
    .X(_2299_));
 sky130_fd_sc_hd__xnor2_1 _6043_ (.A(_2298_),
    .B(_2299_),
    .Y(_2301_));
 sky130_fd_sc_hd__a221o_1 _6044_ (.A1(_2879_),
    .A2(_2296_),
    .B1(_2301_),
    .B2(_2882_),
    .C1(_1025_),
    .X(_2302_));
 sky130_fd_sc_hd__nand2_1 _6045_ (.A(_1502_),
    .B(_1561_),
    .Y(_2303_));
 sky130_fd_sc_hd__or2_1 _6046_ (.A(_1502_),
    .B(_1561_),
    .X(_2304_));
 sky130_fd_sc_hd__a21o_1 _6047_ (.A1(_2303_),
    .A2(_2304_),
    .B1(_1627_),
    .X(_2305_));
 sky130_fd_sc_hd__o211a_1 _6048_ (.A1(_2292_),
    .A2(_2302_),
    .B1(_2305_),
    .C1(_1862_),
    .X(net30));
 sky130_fd_sc_hd__a21oi_1 _6049_ (.A1(_1000_),
    .A2(_1012_),
    .B1(_1980_),
    .Y(_2306_));
 sky130_fd_sc_hd__o21a_1 _6050_ (.A1(_1000_),
    .A2(_1012_),
    .B1(_2306_),
    .X(_2307_));
 sky130_fd_sc_hd__nand2_1 _6051_ (.A(_2811_),
    .B(_2818_),
    .Y(_2308_));
 sky130_fd_sc_hd__or2_1 _6052_ (.A(_2811_),
    .B(_2818_),
    .X(_2309_));
 sky130_fd_sc_hd__and2_1 _6053_ (.A(_2308_),
    .B(_2309_),
    .X(_2311_));
 sky130_fd_sc_hd__nand2_1 _6054_ (.A(_0361_),
    .B(_0365_),
    .Y(_2312_));
 sky130_fd_sc_hd__o21a_1 _6055_ (.A1(_0361_),
    .A2(_0365_),
    .B1(_2885_),
    .X(_2313_));
 sky130_fd_sc_hd__a22o_1 _6056_ (.A1(_2879_),
    .A2(_2311_),
    .B1(_2312_),
    .B2(_2313_),
    .X(_2314_));
 sky130_fd_sc_hd__or2_1 _6057_ (.A(_1469_),
    .B(_1563_),
    .X(_2315_));
 sky130_fd_sc_hd__nand2_1 _6058_ (.A(_1469_),
    .B(_1563_),
    .Y(_2316_));
 sky130_fd_sc_hd__a21o_1 _6059_ (.A1(_2315_),
    .A2(_2316_),
    .B1(_1627_),
    .X(_2317_));
 sky130_fd_sc_hd__o311a_1 _6060_ (.A1(_1025_),
    .A2(_2307_),
    .A3(_2314_),
    .B1(_2317_),
    .C1(_1028_),
    .X(net31));
 sky130_fd_sc_hd__and2b_1 _6061_ (.A_N(_1416_),
    .B(_1564_),
    .X(_2318_));
 sky130_fd_sc_hd__a21oi_1 _6062_ (.A1(_1566_),
    .A2(_2315_),
    .B1(_2318_),
    .Y(_2319_));
 sky130_fd_sc_hd__o21ai_1 _6063_ (.A1(_1416_),
    .A2(_1567_),
    .B1(_1025_),
    .Y(_2321_));
 sky130_fd_sc_hd__xor2_1 _6064_ (.A(_0367_),
    .B(_1796_),
    .X(_2322_));
 sky130_fd_sc_hd__a21bo_1 _6065_ (.A1(_2816_),
    .A2(_2817_),
    .B1_N(_2308_),
    .X(_2323_));
 sky130_fd_sc_hd__xnor2_1 _6066_ (.A(_2323_),
    .B(_2822_),
    .Y(_2324_));
 sky130_fd_sc_hd__o21a_1 _6067_ (.A1(_1000_),
    .A2(_1012_),
    .B1(_1017_),
    .X(_2325_));
 sky130_fd_sc_hd__o21ai_1 _6068_ (.A1(_1009_),
    .A2(_2325_),
    .B1(_2882_),
    .Y(_2326_));
 sky130_fd_sc_hd__a21o_1 _6069_ (.A1(_1009_),
    .A2(_2325_),
    .B1(_2326_),
    .X(_2327_));
 sky130_fd_sc_hd__o211a_1 _6070_ (.A1(_1984_),
    .A2(_2324_),
    .B1(_2327_),
    .C1(_1627_),
    .X(_2328_));
 sky130_fd_sc_hd__o21ai_1 _6071_ (.A1(_2883_),
    .A2(_2322_),
    .B1(_2328_),
    .Y(_2329_));
 sky130_fd_sc_hd__o211a_1 _6072_ (.A1(_2319_),
    .A2(_2321_),
    .B1(_2329_),
    .C1(_1028_),
    .X(net32));
 sky130_fd_sc_hd__or2b_1 _6073_ (.A(_1416_),
    .B_N(_1567_),
    .X(_2331_));
 sky130_fd_sc_hd__xor2_1 _6074_ (.A(_1349_),
    .B(_2331_),
    .X(_2332_));
 sky130_fd_sc_hd__xor2_1 _6075_ (.A(_2617_),
    .B(_2825_),
    .X(_2333_));
 sky130_fd_sc_hd__or3_1 _6076_ (.A(_1020_),
    .B(_1014_),
    .C(_1019_),
    .X(_2334_));
 sky130_fd_sc_hd__a31o_1 _6077_ (.A1(_1021_),
    .A2(_1744_),
    .A3(_2334_),
    .B1(_1024_),
    .X(_2335_));
 sky130_fd_sc_hd__o21ai_1 _6078_ (.A1(_0218_),
    .A2(_0369_),
    .B1(_0149_),
    .Y(_2336_));
 sky130_fd_sc_hd__and3_1 _6079_ (.A(_0370_),
    .B(_2885_),
    .C(_2336_),
    .X(_2337_));
 sky130_fd_sc_hd__a211o_1 _6080_ (.A1(_2879_),
    .A2(_2333_),
    .B1(_2335_),
    .C1(_2337_),
    .X(_2338_));
 sky130_fd_sc_hd__o211a_1 _6081_ (.A1(_1631_),
    .A2(_2332_),
    .B1(_2338_),
    .C1(_1028_),
    .X(net17));
 sky130_fd_sc_hd__or4_1 _6082_ (.A(net1),
    .B(net11),
    .C(net13),
    .D(net12),
    .X(_2339_));
 sky130_fd_sc_hd__buf_2 _6083_ (.A(_2339_),
    .X(_2341_));
 sky130_fd_sc_hd__mux2_1 _6084_ (.A0(net2),
    .A1(_0964_),
    .S(_2341_),
    .X(_2342_));
 sky130_fd_sc_hd__clkbuf_1 _6085_ (.A(_2342_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _6086_ (.A0(net3),
    .A1(_0531_),
    .S(_2341_),
    .X(_2343_));
 sky130_fd_sc_hd__clkbuf_1 _6087_ (.A(_2343_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _6088_ (.A0(net4),
    .A1(_0490_),
    .S(_2341_),
    .X(_2344_));
 sky130_fd_sc_hd__clkbuf_1 _6089_ (.A(_2344_),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _6090_ (.A0(net5),
    .A1(_0533_),
    .S(_2341_),
    .X(_2345_));
 sky130_fd_sc_hd__clkbuf_1 _6091_ (.A(_2345_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _6092_ (.A0(net6),
    .A1(_0581_),
    .S(_2341_),
    .X(_2346_));
 sky130_fd_sc_hd__clkbuf_1 _6093_ (.A(_2346_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _6094_ (.A0(net7),
    .A1(_0573_),
    .S(_2341_),
    .X(_2348_));
 sky130_fd_sc_hd__clkbuf_1 _6095_ (.A(_2348_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _6096_ (.A0(net8),
    .A1(_0697_),
    .S(_2341_),
    .X(_2349_));
 sky130_fd_sc_hd__clkbuf_1 _6097_ (.A(_2349_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _6098_ (.A0(net9),
    .A1(_0698_),
    .S(_2341_),
    .X(_2350_));
 sky130_fd_sc_hd__clkbuf_1 _6099_ (.A(_2350_),
    .X(_0007_));
 sky130_fd_sc_hd__or4b_1 _6100_ (.A(net1),
    .B(net13),
    .C(net12),
    .D_N(net11),
    .X(_2351_));
 sky130_fd_sc_hd__clkbuf_4 _6101_ (.A(_2351_),
    .X(_2352_));
 sky130_fd_sc_hd__mux2_1 _6102_ (.A0(net2),
    .A1(_0899_),
    .S(_2352_),
    .X(_2353_));
 sky130_fd_sc_hd__clkbuf_1 _6103_ (.A(_2353_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _6104_ (.A0(net3),
    .A1(_0720_),
    .S(_2352_),
    .X(_2355_));
 sky130_fd_sc_hd__clkbuf_1 _6105_ (.A(_2355_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _6106_ (.A0(net4),
    .A1(_0421_),
    .S(_2352_),
    .X(_2356_));
 sky130_fd_sc_hd__clkbuf_1 _6107_ (.A(_2356_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _6108_ (.A0(net5),
    .A1(_0506_),
    .S(_2352_),
    .X(_2357_));
 sky130_fd_sc_hd__clkbuf_1 _6109_ (.A(_2357_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _6110_ (.A0(net6),
    .A1(_0671_),
    .S(_2352_),
    .X(_2358_));
 sky130_fd_sc_hd__clkbuf_1 _6111_ (.A(_2358_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _6112_ (.A0(net7),
    .A1(_0684_),
    .S(_2352_),
    .X(_2359_));
 sky130_fd_sc_hd__clkbuf_1 _6113_ (.A(_2359_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _6114_ (.A0(net8),
    .A1(_0546_),
    .S(_2352_),
    .X(_2361_));
 sky130_fd_sc_hd__clkbuf_1 _6115_ (.A(_2361_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _6116_ (.A0(net9),
    .A1(_1585_),
    .S(_2352_),
    .X(_2362_));
 sky130_fd_sc_hd__clkbuf_1 _6117_ (.A(_2362_),
    .X(_0015_));
 sky130_fd_sc_hd__or4b_1 _6118_ (.A(net1),
    .B(net11),
    .C(net13),
    .D_N(net12),
    .X(_2363_));
 sky130_fd_sc_hd__buf_2 _6119_ (.A(_2363_),
    .X(_2364_));
 sky130_fd_sc_hd__mux2_1 _6120_ (.A0(net2),
    .A1(_2550_),
    .S(_2364_),
    .X(_2365_));
 sky130_fd_sc_hd__clkbuf_1 _6121_ (.A(_2365_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _6122_ (.A0(net3),
    .A1(_0883_),
    .S(_2364_),
    .X(_2366_));
 sky130_fd_sc_hd__clkbuf_1 _6123_ (.A(_2366_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _6124_ (.A0(net4),
    .A1(_0971_),
    .S(_2364_),
    .X(_2368_));
 sky130_fd_sc_hd__clkbuf_1 _6125_ (.A(_2368_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _6126_ (.A0(net5),
    .A1(_0916_),
    .S(_2364_),
    .X(_2369_));
 sky130_fd_sc_hd__clkbuf_1 _6127_ (.A(_2369_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _6128_ (.A0(net6),
    .A1(_1915_),
    .S(_2364_),
    .X(_2370_));
 sky130_fd_sc_hd__clkbuf_1 _6129_ (.A(_2370_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _6130_ (.A0(net7),
    .A1(_2445_),
    .S(_2364_),
    .X(_2371_));
 sky130_fd_sc_hd__clkbuf_1 _6131_ (.A(_2371_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _6132_ (.A0(net8),
    .A1(_2858_),
    .S(_2364_),
    .X(_2372_));
 sky130_fd_sc_hd__clkbuf_1 _6133_ (.A(_2372_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _6134_ (.A0(net9),
    .A1(_2859_),
    .S(_2364_),
    .X(_2374_));
 sky130_fd_sc_hd__clkbuf_1 _6135_ (.A(_2374_),
    .X(_0023_));
 sky130_fd_sc_hd__and4bb_4 _6136_ (.A_N(_1028_),
    .B_N(net13),
    .C(net12),
    .D(net11),
    .X(_2375_));
 sky130_fd_sc_hd__mux2_1 _6137_ (.A0(_2717_),
    .A1(net2),
    .S(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__clkbuf_1 _6138_ (.A(_2376_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _6139_ (.A0(_2544_),
    .A1(net3),
    .S(_2375_),
    .X(_2377_));
 sky130_fd_sc_hd__clkbuf_1 _6140_ (.A(_2377_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _6141_ (.A0(_0718_),
    .A1(net4),
    .S(_2375_),
    .X(_2378_));
 sky130_fd_sc_hd__clkbuf_1 _6142_ (.A(_2378_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _6143_ (.A0(_1532_),
    .A1(net5),
    .S(_2375_),
    .X(_2380_));
 sky130_fd_sc_hd__clkbuf_1 _6144_ (.A(_2380_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _6145_ (.A0(_2668_),
    .A1(net6),
    .S(_2375_),
    .X(_2381_));
 sky130_fd_sc_hd__clkbuf_1 _6146_ (.A(_2381_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _6147_ (.A0(_2676_),
    .A1(net7),
    .S(_2375_),
    .X(_2382_));
 sky130_fd_sc_hd__clkbuf_1 _6148_ (.A(_2382_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _6149_ (.A0(_2551_),
    .A1(net8),
    .S(_2375_),
    .X(_2383_));
 sky130_fd_sc_hd__clkbuf_1 _6150_ (.A(_2383_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _6151_ (.A0(_2845_),
    .A1(net9),
    .S(_2375_),
    .X(_2384_));
 sky130_fd_sc_hd__clkbuf_1 _6152_ (.A(_2384_),
    .X(_0031_));
 sky130_fd_sc_hd__or4b_1 _6153_ (.A(net1),
    .B(net11),
    .C(net12),
    .D_N(net13),
    .X(_2386_));
 sky130_fd_sc_hd__buf_2 _6154_ (.A(_2386_),
    .X(_2387_));
 sky130_fd_sc_hd__mux2_1 _6155_ (.A0(net2),
    .A1(_0280_),
    .S(_2387_),
    .X(_2388_));
 sky130_fd_sc_hd__clkbuf_1 _6156_ (.A(_2388_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _6157_ (.A0(net3),
    .A1(_0282_),
    .S(_2387_),
    .X(_2389_));
 sky130_fd_sc_hd__clkbuf_1 _6158_ (.A(_2389_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _6159_ (.A0(net4),
    .A1(_0241_),
    .S(_2387_),
    .X(_2390_));
 sky130_fd_sc_hd__clkbuf_1 _6160_ (.A(_2390_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _6161_ (.A0(net5),
    .A1(_0185_),
    .S(_2387_),
    .X(_2391_));
 sky130_fd_sc_hd__clkbuf_1 _6162_ (.A(_2391_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _6163_ (.A0(net6),
    .A1(_0186_),
    .S(_2387_),
    .X(_2393_));
 sky130_fd_sc_hd__clkbuf_1 _6164_ (.A(_2393_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _6165_ (.A0(net7),
    .A1(_0400_),
    .S(_2387_),
    .X(_2394_));
 sky130_fd_sc_hd__clkbuf_1 _6166_ (.A(_2394_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _6167_ (.A0(net8),
    .A1(_1602_),
    .S(_2387_),
    .X(_2395_));
 sky130_fd_sc_hd__clkbuf_1 _6168_ (.A(_2395_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _6169_ (.A0(net9),
    .A1(_1229_),
    .S(_2387_),
    .X(_2396_));
 sky130_fd_sc_hd__clkbuf_1 _6170_ (.A(_2396_),
    .X(_0039_));
 sky130_fd_sc_hd__and4bb_4 _6171_ (.A_N(_1028_),
    .B_N(net12),
    .C(net13),
    .D(net11),
    .X(_2397_));
 sky130_fd_sc_hd__mux2_1 _6172_ (.A0(_2471_),
    .A1(net2),
    .S(_2397_),
    .X(_2398_));
 sky130_fd_sc_hd__clkbuf_1 _6173_ (.A(_2398_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _6174_ (.A0(_2433_),
    .A1(net3),
    .S(_2397_),
    .X(_2400_));
 sky130_fd_sc_hd__clkbuf_1 _6175_ (.A(_2400_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _6176_ (.A0(_2432_),
    .A1(net4),
    .S(_2397_),
    .X(_2401_));
 sky130_fd_sc_hd__clkbuf_1 _6177_ (.A(_2401_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _6178_ (.A0(_2440_),
    .A1(net5),
    .S(_2397_),
    .X(_2402_));
 sky130_fd_sc_hd__clkbuf_1 _6179_ (.A(_2402_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _6180_ (.A0(_0949_),
    .A1(net6),
    .S(_2397_),
    .X(_2403_));
 sky130_fd_sc_hd__clkbuf_1 _6181_ (.A(_2403_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _6182_ (.A0(_2856_),
    .A1(net7),
    .S(_2397_),
    .X(_2404_));
 sky130_fd_sc_hd__clkbuf_1 _6183_ (.A(_2404_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _6184_ (.A0(_0530_),
    .A1(net8),
    .S(_2397_),
    .X(_2406_));
 sky130_fd_sc_hd__clkbuf_1 _6185_ (.A(_2406_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _6186_ (.A0(_2862_),
    .A1(net9),
    .S(_2397_),
    .X(_2407_));
 sky130_fd_sc_hd__clkbuf_1 _6187_ (.A(_2407_),
    .X(_0047_));
 sky130_fd_sc_hd__and4bb_4 _6188_ (.A_N(net1),
    .B_N(net11),
    .C(net13),
    .D(net12),
    .X(_2408_));
 sky130_fd_sc_hd__mux2_1 _6189_ (.A0(_0342_),
    .A1(net2),
    .S(_2408_),
    .X(_2409_));
 sky130_fd_sc_hd__clkbuf_1 _6190_ (.A(_2409_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _6191_ (.A0(_0293_),
    .A1(net3),
    .S(_2408_),
    .X(_2410_));
 sky130_fd_sc_hd__clkbuf_1 _6192_ (.A(_2410_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _6193_ (.A0(_0294_),
    .A1(net4),
    .S(_2408_),
    .X(_2412_));
 sky130_fd_sc_hd__clkbuf_1 _6194_ (.A(_2412_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _6195_ (.A0(_3002_),
    .A1(net5),
    .S(_2408_),
    .X(_2413_));
 sky130_fd_sc_hd__clkbuf_1 _6196_ (.A(_2413_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _6197_ (.A0(_0229_),
    .A1(net6),
    .S(_2408_),
    .X(_2414_));
 sky130_fd_sc_hd__clkbuf_1 _6198_ (.A(_2414_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _6199_ (.A0(_0378_),
    .A1(net7),
    .S(_2408_),
    .X(_2415_));
 sky130_fd_sc_hd__clkbuf_1 _6200_ (.A(_2415_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _6201_ (.A0(_0388_),
    .A1(net8),
    .S(_2408_),
    .X(_2416_));
 sky130_fd_sc_hd__clkbuf_1 _6202_ (.A(_2416_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _6203_ (.A0(_1029_),
    .A1(net9),
    .S(_2408_),
    .X(_2418_));
 sky130_fd_sc_hd__clkbuf_1 _6204_ (.A(_2418_),
    .X(_0055_));
 sky130_fd_sc_hd__and4b_1 _6205_ (.A_N(net1),
    .B(net11),
    .C(net13),
    .D(net12),
    .X(_2419_));
 sky130_fd_sc_hd__clkbuf_4 _6206_ (.A(_2419_),
    .X(_2420_));
 sky130_fd_sc_hd__mux2_1 _6207_ (.A0(_2778_),
    .A1(net2),
    .S(_2420_),
    .X(_2421_));
 sky130_fd_sc_hd__clkbuf_1 _6208_ (.A(_2421_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _6209_ (.A0(_1235_),
    .A1(net3),
    .S(_2420_),
    .X(_2422_));
 sky130_fd_sc_hd__clkbuf_1 _6210_ (.A(_2422_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _6211_ (.A0(_1806_),
    .A1(net4),
    .S(_2420_),
    .X(_2423_));
 sky130_fd_sc_hd__clkbuf_1 _6212_ (.A(_2423_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _6213_ (.A0(_2347_),
    .A1(net5),
    .S(_2420_),
    .X(_2425_));
 sky130_fd_sc_hd__clkbuf_1 _6214_ (.A(_2425_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _6215_ (.A0(_2630_),
    .A1(net6),
    .S(_2420_),
    .X(_2426_));
 sky130_fd_sc_hd__clkbuf_1 _6216_ (.A(_2426_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _6217_ (.A0(_1521_),
    .A1(net7),
    .S(_2420_),
    .X(_2427_));
 sky130_fd_sc_hd__clkbuf_1 _6218_ (.A(_2427_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _6219_ (.A0(_2833_),
    .A1(net8),
    .S(_2420_),
    .X(_2428_));
 sky130_fd_sc_hd__clkbuf_1 _6220_ (.A(_2428_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _6221_ (.A0(_0696_),
    .A1(net9),
    .S(_2420_),
    .X(_2429_));
 sky130_fd_sc_hd__clkbuf_1 _6222_ (.A(_2429_),
    .X(_0063_));
 sky130_fd_sc_hd__dfrtp_1 _6223_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0000_),
    .RESET_B(net39),
    .Q(\A[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _6224_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0001_),
    .RESET_B(net39),
    .Q(\A[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _6225_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0002_),
    .RESET_B(net39),
    .Q(\A[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _6226_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0003_),
    .RESET_B(net39),
    .Q(\A[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _6227_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0004_),
    .RESET_B(net39),
    .Q(\A[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6228_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0005_),
    .RESET_B(net39),
    .Q(\A[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6229_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0006_),
    .RESET_B(net39),
    .Q(\A[0][6] ));
 sky130_fd_sc_hd__dfrtp_4 _6230_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0007_),
    .RESET_B(net39),
    .Q(\A[0][7] ));
 sky130_fd_sc_hd__dfrtp_4 _6231_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0008_),
    .RESET_B(net35),
    .Q(\A[1][0] ));
 sky130_fd_sc_hd__dfrtp_1 _6232_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0009_),
    .RESET_B(net33),
    .Q(\A[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _6233_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0010_),
    .RESET_B(net35),
    .Q(\A[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _6234_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0011_),
    .RESET_B(net35),
    .Q(\A[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _6235_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0012_),
    .RESET_B(net35),
    .Q(\A[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6236_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0013_),
    .RESET_B(net35),
    .Q(\A[1][5] ));
 sky130_fd_sc_hd__dfrtp_1 _6237_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0014_),
    .RESET_B(net35),
    .Q(\A[1][6] ));
 sky130_fd_sc_hd__dfrtp_4 _6238_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0015_),
    .RESET_B(net36),
    .Q(\A[1][7] ));
 sky130_fd_sc_hd__dfrtp_1 _6239_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0016_),
    .RESET_B(net37),
    .Q(\A[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _6240_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0017_),
    .RESET_B(net37),
    .Q(\A[2][1] ));
 sky130_fd_sc_hd__dfrtp_1 _6241_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0018_),
    .RESET_B(net37),
    .Q(\A[2][2] ));
 sky130_fd_sc_hd__dfrtp_1 _6242_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0019_),
    .RESET_B(net37),
    .Q(\A[2][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6243_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0020_),
    .RESET_B(net37),
    .Q(\A[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6244_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0021_),
    .RESET_B(net37),
    .Q(\A[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _6245_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0022_),
    .RESET_B(net37),
    .Q(\A[2][6] ));
 sky130_fd_sc_hd__dfrtp_4 _6246_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0023_),
    .RESET_B(net38),
    .Q(\A[2][7] ));
 sky130_fd_sc_hd__dfrtp_1 _6247_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0024_),
    .RESET_B(net33),
    .Q(\A[3][0] ));
 sky130_fd_sc_hd__dfrtp_1 _6248_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0025_),
    .RESET_B(net33),
    .Q(\A[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _6249_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0026_),
    .RESET_B(net33),
    .Q(\A[3][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6250_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0027_),
    .RESET_B(net33),
    .Q(\A[3][3] ));
 sky130_fd_sc_hd__dfrtp_1 _6251_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0028_),
    .RESET_B(net33),
    .Q(\A[3][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6252_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0029_),
    .RESET_B(net34),
    .Q(\A[3][5] ));
 sky130_fd_sc_hd__dfrtp_1 _6253_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0030_),
    .RESET_B(net34),
    .Q(\A[3][6] ));
 sky130_fd_sc_hd__dfrtp_4 _6254_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0031_),
    .RESET_B(net36),
    .Q(\A[3][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6255_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0032_),
    .RESET_B(net38),
    .Q(\B[0][0] ));
 sky130_fd_sc_hd__dfrtp_4 _6256_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0033_),
    .RESET_B(net38),
    .Q(\B[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _6257_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0034_),
    .RESET_B(net38),
    .Q(\B[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _6258_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0035_),
    .RESET_B(net38),
    .Q(\B[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _6259_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0036_),
    .RESET_B(net38),
    .Q(\B[0][4] ));
 sky130_fd_sc_hd__dfrtp_4 _6260_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0037_),
    .RESET_B(net39),
    .Q(\B[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6261_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0038_),
    .RESET_B(net37),
    .Q(\B[0][6] ));
 sky130_fd_sc_hd__dfrtp_4 _6262_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0039_),
    .RESET_B(net37),
    .Q(\B[0][7] ));
 sky130_fd_sc_hd__dfrtp_1 _6263_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0040_),
    .RESET_B(net37),
    .Q(\B[1][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6264_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0041_),
    .RESET_B(net40),
    .Q(\B[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _6265_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0042_),
    .RESET_B(net39),
    .Q(\B[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _6266_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0043_),
    .RESET_B(net40),
    .Q(\B[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _6267_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0044_),
    .RESET_B(net40),
    .Q(\B[1][4] ));
 sky130_fd_sc_hd__dfrtp_4 _6268_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0045_),
    .RESET_B(net40),
    .Q(\B[1][5] ));
 sky130_fd_sc_hd__dfrtp_4 _6269_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0046_),
    .RESET_B(net40),
    .Q(\B[1][6] ));
 sky130_fd_sc_hd__dfrtp_4 _6270_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0047_),
    .RESET_B(net40),
    .Q(\B[1][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6271_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0048_),
    .RESET_B(net40),
    .Q(\B[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _6272_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0049_),
    .RESET_B(net33),
    .Q(\B[2][1] ));
 sky130_fd_sc_hd__dfrtp_4 _6273_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0050_),
    .RESET_B(net34),
    .Q(\B[2][2] ));
 sky130_fd_sc_hd__dfrtp_4 _6274_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0051_),
    .RESET_B(net34),
    .Q(\B[2][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6275_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0052_),
    .RESET_B(net34),
    .Q(\B[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _6276_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0053_),
    .RESET_B(net34),
    .Q(\B[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _6277_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0054_),
    .RESET_B(net34),
    .Q(\B[2][6] ));
 sky130_fd_sc_hd__dfrtp_4 _6278_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0055_),
    .RESET_B(net34),
    .Q(\B[2][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6279_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0056_),
    .RESET_B(net36),
    .Q(\B[3][0] ));
 sky130_fd_sc_hd__dfrtp_1 _6280_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0057_),
    .RESET_B(net33),
    .Q(\B[3][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6281_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0058_),
    .RESET_B(net35),
    .Q(\B[3][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6282_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0059_),
    .RESET_B(net33),
    .Q(\B[3][3] ));
 sky130_fd_sc_hd__dfrtp_4 _6283_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0060_),
    .RESET_B(net33),
    .Q(\B[3][4] ));
 sky130_fd_sc_hd__dfrtp_4 _6284_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0061_),
    .RESET_B(net35),
    .Q(\B[3][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6285_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0062_),
    .RESET_B(net35),
    .Q(\B[3][6] ));
 sky130_fd_sc_hd__dfrtp_4 _6286_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0063_),
    .RESET_B(net36),
    .Q(\B[3][7] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(execute),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input2 (.A(input_val[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(input_val[1]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(input_val[2]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(input_val[3]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(input_val[4]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(input_val[5]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(input_val[6]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(input_val[7]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input10 (.A(reset),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(sel_in[0]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(sel_in[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(sel_in[2]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(sel_out[0]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(sel_out[1]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(out[0]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(out[10]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(out[11]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(out[12]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(out[13]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(out[14]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(out[15]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(out[16]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(out[1]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(out[2]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(out[3]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(out[4]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(out[5]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(out[6]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(out[7]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(out[8]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(out[9]));
 sky130_fd_sc_hd__clkbuf_4 fanout33 (.A(net34),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 fanout36 (.A(net10),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 fanout37 (.A(net40),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(net40),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__buf_4 fanout40 (.A(net10),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\B[1][2] ),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\B[3][1] ),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\A[2][4] ),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\B[1][1] ),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\B[3][5] ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\A[0][4] ),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\A[2][1] ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\B[2][6] ),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\A[3][2] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\A[2][5] ),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\A[3][4] ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\A[0][3] ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\A[0][2] ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\B[0][2] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\A[3][5] ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\A[0][6] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\A[2][3] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\A[2][2] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\B[0][3] ),
    .X(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__C (.DIODE(\A[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__B (.DIODE(\A[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A2 (.DIODE(\A[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__A (.DIODE(\A[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__A1_N (.DIODE(\A[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A2 (.DIODE(\A[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__A (.DIODE(\A[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__C (.DIODE(\A[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__B (.DIODE(\A[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__B (.DIODE(\A[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A (.DIODE(\A[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__A (.DIODE(\A[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A1 (.DIODE(\A[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__A1 (.DIODE(\A[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__A1 (.DIODE(\A[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__A1 (.DIODE(\A[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__A (.DIODE(\A[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__A1 (.DIODE(\A[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__A (.DIODE(\A[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__A (.DIODE(\A[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A1 (.DIODE(\A[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A1 (.DIODE(\A[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A (.DIODE(\A[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__A (.DIODE(\A[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__A1 (.DIODE(\A[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__A (.DIODE(\A[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3271__A (.DIODE(\A[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__D (.DIODE(\A[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__B1 (.DIODE(\A[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__C (.DIODE(\A[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A2 (.DIODE(\A[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__B (.DIODE(\A[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__D (.DIODE(\A[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__C (.DIODE(\A[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__A2 (.DIODE(\A[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__A (.DIODE(\A[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A1 (.DIODE(\A[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__A (.DIODE(\A[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A (.DIODE(\A[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A1 (.DIODE(\A[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__A1 (.DIODE(\A[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__A1 (.DIODE(\A[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__A (.DIODE(\A[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__A1 (.DIODE(\A[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__A (.DIODE(\A[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A (.DIODE(\B[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__B (.DIODE(\B[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__B (.DIODE(\B[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__A1 (.DIODE(\B[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__C (.DIODE(\B[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__D (.DIODE(\B[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__C (.DIODE(\B[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__A (.DIODE(\B[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A (.DIODE(\B[0][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A (.DIODE(\B[0][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A (.DIODE(\B[0][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A (.DIODE(\B[0][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A1 (.DIODE(\B[0][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__A (.DIODE(\B[0][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__B (.DIODE(\B[0][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__B (.DIODE(\B[0][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__B (.DIODE(\B[0][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__B (.DIODE(\B[0][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A1 (.DIODE(\B[0][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__B (.DIODE(\B[0][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A (.DIODE(\B[0][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__B (.DIODE(\B[0][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A1 (.DIODE(\B[0][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__A (.DIODE(\B[1][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__C (.DIODE(\B[1][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__A (.DIODE(\B[1][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__A (.DIODE(\B[1][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__A (.DIODE(\B[1][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__A (.DIODE(\B[1][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__A (.DIODE(\B[1][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__A (.DIODE(\B[1][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__B2 (.DIODE(\B[1][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A (.DIODE(\B[1][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__A (.DIODE(\B[1][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__A (.DIODE(\B[1][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__B2 (.DIODE(\B[1][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__A (.DIODE(\B[1][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__B (.DIODE(\B[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__A1 (.DIODE(\B[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__B (.DIODE(\B[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3294__B (.DIODE(\B[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__B (.DIODE(\B[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__A1 (.DIODE(\B[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__B (.DIODE(\B[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3220__A (.DIODE(\B[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__B (.DIODE(\B[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__A1 (.DIODE(\B[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__A (.DIODE(\B[2][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__A2 (.DIODE(\B[2][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__B (.DIODE(\B[2][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__C (.DIODE(\B[2][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__D (.DIODE(\B[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__A2 (.DIODE(\B[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__B (.DIODE(\B[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A (.DIODE(\B[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__B1 (.DIODE(\B[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__B (.DIODE(\B[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A (.DIODE(\B[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__A (.DIODE(\B[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__B (.DIODE(\B[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__D (.DIODE(\B[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__C (.DIODE(\B[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A2 (.DIODE(\B[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__D (.DIODE(\B[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__C (.DIODE(\B[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__A (.DIODE(\B[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A (.DIODE(\B[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A (.DIODE(\B[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A (.DIODE(\B[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A (.DIODE(\B[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__A2 (.DIODE(\B[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__B (.DIODE(\B[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3120__A2 (.DIODE(\B[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3113__A (.DIODE(\B[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__C (.DIODE(\B[3][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__D (.DIODE(\B[3][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__B (.DIODE(\B[3][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3177__C (.DIODE(\B[3][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__A (.DIODE(\B[3][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3142__A (.DIODE(\B[3][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__B (.DIODE(\B[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__B (.DIODE(\B[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3174__B (.DIODE(\B[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3151__A (.DIODE(\B[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__B (.DIODE(\B[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__D (.DIODE(\B[3][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__D (.DIODE(\B[3][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__D (.DIODE(\B[3][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__A (.DIODE(\B[3][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__D (.DIODE(\B[3][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__A (.DIODE(\B[3][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold5_A (.DIODE(\B[3][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__A (.DIODE(\B[3][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__A (.DIODE(\B[3][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__A (.DIODE(\B[3][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__A (.DIODE(\B[3][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__A1 (.DIODE(\B[3][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__A (.DIODE(\B[3][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__A (.DIODE(\B[3][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__A (.DIODE(\B[3][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3161__A (.DIODE(\B[3][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__A (.DIODE(\B[3][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__A (.DIODE(\B[3][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__A (.DIODE(\B[3][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A (.DIODE(\B[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__A (.DIODE(\B[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A (.DIODE(\B[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__A (.DIODE(\B[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3235__A (.DIODE(\B[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__A (.DIODE(\B[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__B (.DIODE(_0071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A2 (.DIODE(_0071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__B1 (.DIODE(_0072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A1 (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__A1 (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__A (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__A1 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__A (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A2 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__B (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__A (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__A (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__A1 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__A1 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A2 (.DIODE(_0085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__B (.DIODE(_0085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__B1 (.DIODE(_0085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A2 (.DIODE(_0085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__D (.DIODE(_0085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__B (.DIODE(_0085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A (.DIODE(_0085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A2 (.DIODE(_0085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__B (.DIODE(_0085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A2 (.DIODE(_0085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__B1 (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__B (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__B (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__A2 (.DIODE(_0140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__C (.DIODE(_0140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A2 (.DIODE(_0140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__A1 (.DIODE(_0141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__A (.DIODE(_0141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__B1_N (.DIODE(_0141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A2 (.DIODE(_0148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__A2 (.DIODE(_0148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__B (.DIODE(_0148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__B1 (.DIODE(_0150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__A (.DIODE(_0150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A (.DIODE(_0151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__A (.DIODE(_0151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__C (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__C (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__A2 (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__B (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__A2 (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__B (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__A1 (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__A2 (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__C (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__C (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__D (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__D (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__B1 (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__D (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__B2 (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__B1 (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__B1 (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__D (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__A (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__D (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__A (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__B1 (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__B (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__B (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__A (.DIODE(_0159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A1 (.DIODE(_0159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A1 (.DIODE(_0159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A (.DIODE(_0159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A1 (.DIODE(_0159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__A (.DIODE(_0159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__A (.DIODE(_0159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A1 (.DIODE(_0159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__A (.DIODE(_0159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__A1 (.DIODE(_0159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__D (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__D (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__B2 (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__B (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__B1 (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__B1 (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__D (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__B2 (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__D (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__B2 (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__B1 (.DIODE(_0181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__A1 (.DIODE(_0181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__C1 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__A2 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__A1 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__B (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__C (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__C (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__B (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__B (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__B (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__A2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A1 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__B1 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__B1 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__D (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__B1 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__D (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__B (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__D (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__B1 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__B1 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__A1 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__A (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__A (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__A2 (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__C (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__C (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__D (.DIODE(_0220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__C (.DIODE(_0220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__B (.DIODE(_0220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__D (.DIODE(_0220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__C (.DIODE(_0220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A2 (.DIODE(_0220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__B1 (.DIODE(_0220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__B1 (.DIODE(_0220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__C (.DIODE(_0220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__A2 (.DIODE(_0220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__B (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__C (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__A2 (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__B (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__A2 (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__A2 (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__B (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__B2 (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__A0 (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__B (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A2 (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__B (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__B2 (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__B2 (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__B1 (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__D (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__B (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__B (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__A1 (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__B (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A2 (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__B (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__B1 (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__A (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__B (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__B (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A2 (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__B1 (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__B1 (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__A1 (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__C (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A1 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__A (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__A (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__A (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__A (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__A (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__A1 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__A (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__A1 (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__B (.DIODE(_0275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__A2 (.DIODE(_0275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__A (.DIODE(_0278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__A (.DIODE(_0278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A (.DIODE(_0279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__B2 (.DIODE(_0279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__B2 (.DIODE(_0279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A (.DIODE(_0279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__B2 (.DIODE(_0279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__A2 (.DIODE(_0279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__C (.DIODE(_0279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__A2 (.DIODE(_0279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__A2 (.DIODE(_0279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__A (.DIODE(_0279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A1 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__A1 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A1 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A1 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__C (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__A (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__B2 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__A (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__A1 (.DIODE(_0282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__B1 (.DIODE(_0282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__D (.DIODE(_0282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__B (.DIODE(_0282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A2 (.DIODE(_0282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__B1 (.DIODE(_0282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__B1 (.DIODE(_0282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__D (.DIODE(_0282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__A2 (.DIODE(_0282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__C (.DIODE(_0282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__A0 (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__B (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A2 (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__C (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A1 (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__B2 (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__B2 (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__B (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__A1 (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__B (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__A0 (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__B1 (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__D (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__B1 (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A2 (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A1 (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__B (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__B1 (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__B1 (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__D (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__A0 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__B1 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__B2 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__C (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A1 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__B (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__A1 (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A1 (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__B1 (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__A0 (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__A (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__A1 (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A1 (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A1 (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__A1 (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__A (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__A1 (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__A (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__B1_N (.DIODE(_0381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__B (.DIODE(_0381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__A (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__A (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__A0 (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__B (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__B (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__B2 (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__B (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__B1 (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A1 (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__A (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__A1 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A1 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A1 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A1 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__A1_N (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__A1 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__A1 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__A1 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A2 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__B2 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__B (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__A1 (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__B (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__B (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A1_N (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__B (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__A2 (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A2 (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__B (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__B (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A2 (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__B2 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__B (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__B2 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__B (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B2 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__A (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__A (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__B2 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__A (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__A (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A1 (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__A (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__A2 (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__A (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__B2 (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__A (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__A (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__B (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__C (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A1 (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A1 (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__A (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__A (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A1 (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__A (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__A (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__A (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A2 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__B (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__D (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__B (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__B (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__B (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__C (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__D (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__A1 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__B1 (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__B (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__B (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__B2 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__A2 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__B1 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__C (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__B (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__A (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__C (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__A2 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A1 (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A1 (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__B1 (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__B (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__B2 (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A2_N (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__A2 (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__D (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__D (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__B1 (.DIODE(_0490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__B1 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__B (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A2 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__B (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A2 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__C (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__B1 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__A (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__B (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__B (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A2 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A1 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__B (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__B2 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__A (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__A (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__A (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__A1 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__A (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__A1 (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A2 (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__B (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__B (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__B (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__B (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__A2 (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__B (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__A2 (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__B (.DIODE(_0506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__A0 (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__C (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__C (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A2 (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A2 (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__B (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__B (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__B (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__A (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__A1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A2 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__C (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__A2_N (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__D (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__A2 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__C (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__A1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__C (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__A1 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__B1 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__B2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__A1 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__B (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__B (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__A2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__B1 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__A1 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__A1 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__C (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A1 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__C (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__B2 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__B2 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__B2 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__B2 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__B (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__A (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__A (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__A (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__A (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__B (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__B (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__B2 (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__B2 (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__B (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__B2 (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__B (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__B (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__A (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__B2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__A (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__B2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__A (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A1 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__A1 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__A (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A1 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__B (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__A (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__B (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A2 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A2 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__B (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A1 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__A (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__A1 (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__B1 (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__C (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__B1 (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__C (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__B (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__A2 (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__B (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__B2 (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__B (.DIODE(_0581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__B (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A2 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__B (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A2 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__B (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__A2 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__B (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__A2 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__B (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__B (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__B (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__B (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__A (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__A (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__A (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A1 (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__A (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__A (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3104__A (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__A1 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A1 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__A2 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__B (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__B (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A1 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__A1 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__A (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A2 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__B (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__A2 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__A1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__A1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__A1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__A (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A0 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A2 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A2 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A2 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A2 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__A (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__A1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__A1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__A1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__B (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__C (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A2 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__A (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A2 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__A (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A1 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__B1 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__B1 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A_N (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__B2 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__B2 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__B1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__B1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A2 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__B (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A2 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__C (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__B1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__B (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__A2 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3107__A (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__A2 (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A2 (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__B (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__A0 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__B (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__B (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__B (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A2 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A2 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__B (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__B (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__A2 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__B (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__B (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A1_N (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__C (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__B1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__C (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A2 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__B (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__B (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__B (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__A (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A2 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__B (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__B (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A2 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A2 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__B (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__A2 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__B (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__B2 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__B (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__A2 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__C (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__A1 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__A (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__A2 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__B2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__B2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3294__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__B2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__B2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3109__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__B1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__B (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__B (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__B (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__B (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__A1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A2 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__A (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__A (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__A1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__A1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__A (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__C (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A1 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__B (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__B (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__B (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__A (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__B2 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__B (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__A (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__B (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A1 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__B (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__C (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A1 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__B (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__C (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__A2 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3112__A (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__B (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__B2 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__B1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__D (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__B (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__B2 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__C (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__A2 (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__B (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B1 (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__D (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A2 (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__B (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__B1 (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__B (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__D (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__A2 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__C (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A2 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__A1 (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__A (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__B1_N (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__B (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__B2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__A (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__A (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__A (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__A (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__A (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3120__A1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__A (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__B2 (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A1_N (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__B (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__B (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__B2 (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__A (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__A (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__A (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__B2 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__C (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A2 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__B (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__B (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__A (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__C (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__D (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__B1 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__B (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__B1 (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__B (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__A (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__B2 (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__B1 (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A1 (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__B (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__B1 (.DIODE(_0866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__D (.DIODE(_0866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__A (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__A1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__A (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__C (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__A1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__B1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__D (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__A1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__B (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A2 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__C (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__A1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__A2 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__B (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__A1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__B2 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__B2 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__D (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__A2 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__B (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__A2 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__A (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__B (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__A1 (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__B (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__B (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__A2 (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__B1 (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3303__B (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__B (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__A2 (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__B1 (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__A1 (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__B1 (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__A1 (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__A2 (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__C (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__A2 (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__A1 (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__A2 (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__C (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__C (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__C (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__A1 (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__A2 (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__D (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__D (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__B2 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__D (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__B1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__B1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__D (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__B2 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__D (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__A (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A0 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__B1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__D (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__B1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__B1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__C (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__B1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__B1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__D (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__B1 (.DIODE(_0949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__A1 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__A2 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A1 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__B (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__B2 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A2 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__B2 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__A (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__B2 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__B1 (.DIODE(_0966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__C (.DIODE(_0966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__A1 (.DIODE(_0971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__B (.DIODE(_0971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__B1 (.DIODE(_0971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A2 (.DIODE(_0971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__B (.DIODE(_0971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__A2 (.DIODE(_0971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__D (.DIODE(_0971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__B1 (.DIODE(_0971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__A2 (.DIODE(_0971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__B2 (.DIODE(_0971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__D (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__B1 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__A1 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__C (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__D (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__B2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__A1 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__C (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__A (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__C (.DIODE(_1015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__A2 (.DIODE(_1015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__C (.DIODE(_1015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__A2 (.DIODE(_1015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__A (.DIODE(_1015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__A2 (.DIODE(_1015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__B (.DIODE(_1015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__A2 (.DIODE(_1015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__B (.DIODE(_1015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__C (.DIODE(_1015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__B1 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6026__A (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__B1 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__B1 (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__A (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__B1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__C1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__A (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__C1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__C1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__B1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__B1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__C1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__B1 (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__D (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__B1 (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__B1 (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__B1 (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__D (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__B (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__D (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__B1 (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__D (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__A_N (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__A_N (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__C1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__C1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__C1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__A (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__C1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__C1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__B1 (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__A0 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A2 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__A1 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__A1 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__A1 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A1 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__A1 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A1 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__A1 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__B1 (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3171__A (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__B2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__A (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__A (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__B (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__C (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__A2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3177__B (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__C (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__A2 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__A1 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__B1 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__B1 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__D (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__D (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__A2 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3176__B1 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__B1 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__D (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__B1 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__B (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__B2 (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__A2 (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__A2 (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__C (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__B2 (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__B (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__B2 (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3176__A2 (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__C (.DIODE(_1136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__B_N (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__D (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__B (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__B1 (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__B (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4310__A (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__A2 (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3257__A (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__B1 (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__B (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__A (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__A (.DIODE(_1209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__B (.DIODE(_1209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__B (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__B1 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__B2 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__A (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3255__B (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__C (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__A2 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__C (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__B1 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__B (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__A1 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__B (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__D (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__C1 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__C1 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__A (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__B (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__B2 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A1 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A0 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__B (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A2 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__C (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__A1 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__B (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A2 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__C (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A1 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__A2 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__A2 (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__D (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__B (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__C (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__B1 (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__A2 (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__C (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__A1 (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__A (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__D (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__A (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__A1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__B (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__B (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__A1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__A1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__A (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__A1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__A1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__A (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__A1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__D (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__D (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__B2 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__B2 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__D (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__B2 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__B1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__D (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__D (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__B2 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A1 (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__C (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A2 (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__B (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__A (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__A (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A1 (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__B1 (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__C1 (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A2 (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__B2 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__B1 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A1 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__B1 (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__D (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__D (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A_N (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__B (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__B1 (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__B1 (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A1 (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__C (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__B2 (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__D (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A2 (.DIODE(_1450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__C1 (.DIODE(_1450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A2 (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__B (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A1 (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A1 (.DIODE(_1481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A (.DIODE(_1481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__B1_N (.DIODE(_1481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__C (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__A0 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A2 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A2 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__A (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__A2 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__A (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__A1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__B1 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__C (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A0 (.DIODE(_1532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__A2 (.DIODE(_1532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__B (.DIODE(_1532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__B (.DIODE(_1532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__B (.DIODE(_1532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A2 (.DIODE(_1532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__B (.DIODE(_1532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3235__B (.DIODE(_1532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__B (.DIODE(_1532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__B1 (.DIODE(_1532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__B2 (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__D (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__B2 (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__B1 (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__B (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__B2 (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__A (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__A1 (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__B1 (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__B2 (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__B_N (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__A2 (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__C_N (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__A (.DIODE(_1587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__A (.DIODE(_1587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__A (.DIODE(_1587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__A (.DIODE(_1587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__A (.DIODE(_1587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__A (.DIODE(_1587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3409__A (.DIODE(_1587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3255__A (.DIODE(_1587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__A (.DIODE(_1587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3189__A (.DIODE(_1587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A1 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__A (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__B (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__A1 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A1 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__A (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__A (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__A (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__B (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A1 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__B (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__C (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__B1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__B (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__B (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__B1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__A (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__A (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3189__B (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__C1 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__B1 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__B1 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__C1 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__C1 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__B1 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__A (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__B1 (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__C1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__A1 (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__A1 (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__A1 (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__A1 (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__C1 (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__A1 (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A1 (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A1 (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A1 (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A1 (.DIODE(_1631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A2 (.DIODE(_1688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__B1 (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__A2 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__A2 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A2 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__A2 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__B (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A2 (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A2 (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__B1 (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__B1 (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__A1 (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__B (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__C (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__B1 (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A (.DIODE(_1792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__A1 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A1 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__B (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__B (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__A0 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__B1 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__D (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__B1 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__A2 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__B (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__B1 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__D (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__B1 (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__B (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__A2 (.DIODE(_1856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A2 (.DIODE(_1856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__B (.DIODE(_1856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__A2 (.DIODE(_1856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__B (.DIODE(_1856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__C1 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__C1 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__C1 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__C1 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__C1 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__C1 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__C1 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__C1 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__C1 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__C1 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A2 (.DIODE(_1901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A1_N (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__A (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__A1 (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__A (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__A (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3303__A (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__A (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__A1 (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__A1 (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__A1 (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__B1 (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__B (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__B2 (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__B (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3294__D (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__B (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__B1 (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__C (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__A2 (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__B (.DIODE(_1959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__B (.DIODE(_1959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__A (.DIODE(_1959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__A1 (.DIODE(_1959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__B (.DIODE(_1959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__A1 (.DIODE(_1959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__B (.DIODE(_1959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A (.DIODE(_1959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__A (.DIODE(_1959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__A1 (.DIODE(_1959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__B (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__A1 (.DIODE(_1984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__A2 (.DIODE(_1984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__B1 (.DIODE(_1984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__B1 (.DIODE(_1984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__B1 (.DIODE(_1984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A1 (.DIODE(_1984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A2 (.DIODE(_2047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A1 (.DIODE(_2116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A1 (.DIODE(_2116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__A1 (.DIODE(_2116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A (.DIODE(_2116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A1 (.DIODE(_2118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__C1 (.DIODE(_2118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A2 (.DIODE(_2139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A3 (.DIODE(_2140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A3 (.DIODE(_2179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__B (.DIODE(_2179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__A (.DIODE(_2181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A (.DIODE(_2181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__B1 (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__B (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A1 (.DIODE(_2189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A2 (.DIODE(_2191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A2 (.DIODE(_2197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__B (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__B (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__B (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__B2 (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__A (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__A (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__B (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__B2 (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__A (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__A1 (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__B1 (.DIODE(_2305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__B1 (.DIODE(_2317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__A1 (.DIODE(_2319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__A2 (.DIODE(_2333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A0 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__A2_N (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A2 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__B (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__B (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__B (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__A2_N (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__B (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__D (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__B (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__S (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__S (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__S (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__S (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__S (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__S (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__S (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__S (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__S (.DIODE(_2375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__S (.DIODE(_2375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__S (.DIODE(_2375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__S (.DIODE(_2375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__S (.DIODE(_2375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__S (.DIODE(_2375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__S (.DIODE(_2375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__S (.DIODE(_2375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__A1 (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__B (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__B2 (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__B2 (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__A (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__A (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__A (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__A (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__B (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__A1 (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__A (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__A1 (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__B (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__B2 (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__B2 (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__B (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__A (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3274__A (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__A (.DIODE(_2405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__S (.DIODE(_2408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__S (.DIODE(_2408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__S (.DIODE(_2408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__S (.DIODE(_2408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__S (.DIODE(_2408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__S (.DIODE(_2408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__S (.DIODE(_2408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__S (.DIODE(_2408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__S (.DIODE(_2420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__S (.DIODE(_2420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__S (.DIODE(_2420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__S (.DIODE(_2420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__S (.DIODE(_2420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__S (.DIODE(_2420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__S (.DIODE(_2420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__S (.DIODE(_2420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__B (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__A (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__A (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__A (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__A (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__A1 (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__A (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__A (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__A (.DIODE(_2431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A0 (.DIODE(_2432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__B (.DIODE(_2432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__A2 (.DIODE(_2432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__A (.DIODE(_2432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__A2 (.DIODE(_2432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__B (.DIODE(_2432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__B (.DIODE(_2432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A2 (.DIODE(_2432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__B1 (.DIODE(_2432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__B (.DIODE(_2432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A0 (.DIODE(_2433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__B1 (.DIODE(_2433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__D (.DIODE(_2433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__B1 (.DIODE(_2433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__B (.DIODE(_2433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__B1 (.DIODE(_2433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__D (.DIODE(_2433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__D (.DIODE(_2433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__A2 (.DIODE(_2433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3274__B (.DIODE(_2433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__A1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__C (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__D (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__A2 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A2 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__C (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__B (.DIODE(_2438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__A (.DIODE(_2438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__B (.DIODE(_2438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__B1 (.DIODE(_2438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__B (.DIODE(_2438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__B (.DIODE(_2438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__A (.DIODE(_2438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__A (.DIODE(_2438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__B (.DIODE(_2438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__D (.DIODE(_2438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__A0 (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__B (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__A2 (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__C (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__B2 (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__A1 (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__A2 (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__B (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__A2 (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__B (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__A1 (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__A2 (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__A2 (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__A2 (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__A (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__A2 (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__B2 (.DIODE(_2468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__B (.DIODE(_2468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__A2 (.DIODE(_2468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__A2 (.DIODE(_2468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__C (.DIODE(_2468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__A2 (.DIODE(_2468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__A (.DIODE(_2468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__B2 (.DIODE(_2468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__A2 (.DIODE(_2468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__A2 (.DIODE(_2468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__A (.DIODE(_2470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__B2 (.DIODE(_2470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__B2 (.DIODE(_2470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__A (.DIODE(_2470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__C (.DIODE(_2470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__B2 (.DIODE(_2470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__B2 (.DIODE(_2470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__A2 (.DIODE(_2470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__C (.DIODE(_2470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3311__A (.DIODE(_2470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__A0 (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A1 (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A2 (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__C (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__A1 (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__B (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__A (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A1 (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__C (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__A2 (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__A1 (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__B (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__D (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__C (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__C (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__A1 (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__A1 (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__B1 (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__D (.DIODE(_2496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__B (.DIODE(_2536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__A2 (.DIODE(_2536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__B1 (.DIODE(_2537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__A0 (.DIODE(_2544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__A2 (.DIODE(_2544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__A2 (.DIODE(_2544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__B (.DIODE(_2544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__A2 (.DIODE(_2544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__A2 (.DIODE(_2544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A1 (.DIODE(_2544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__B (.DIODE(_2544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__B (.DIODE(_2544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A2 (.DIODE(_2544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A (.DIODE(_2545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__A1 (.DIODE(_2545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__B (.DIODE(_2545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__A1 (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A2 (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A2 (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__C (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__A1 (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__A (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__B (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__B2 (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__A (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__A2 (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__A0 (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A1 (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__C (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__B (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__B1 (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__D (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__B1 (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__A2 (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__B (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__B2 (.DIODE(_2551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__B1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__B (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__B (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A2 (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__C (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__A2 (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A1 (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__A (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__B1_N (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A0 (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__B (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__B (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__B (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A2 (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__B (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__A2 (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__B2 (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__B (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__B (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__A1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__A1 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A0 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__A2 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__B (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__A2 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__B (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A2 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__B (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A2 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__A2 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__B (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__B (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__B1 (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__B (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A (.DIODE(_2675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__A0 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A1 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__A2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__B (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__B (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__C (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A1 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__B (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A1 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__A (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__A (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__A1 (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__A (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__C (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__A2 (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__C (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A0 (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__B1 (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__B1 (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__A (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__D (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__A2 (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__B (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__A2 (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__B (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__A (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A1 (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__B (.DIODE(_2730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A2 (.DIODE(_2730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__A (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__A (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__A0 (.DIODE(_2778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__B2 (.DIODE(_2778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__B1 (.DIODE(_2778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__D (.DIODE(_2778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A1 (.DIODE(_2778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A (.DIODE(_2778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__D (.DIODE(_2778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__A1 (.DIODE(_2778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__A (.DIODE(_2778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A1 (.DIODE(_2778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A0 (.DIODE(_2833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__B (.DIODE(_2833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__B (.DIODE(_2833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__B2 (.DIODE(_2833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__B1 (.DIODE(_2833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__B (.DIODE(_2833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__B (.DIODE(_2833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__A1 (.DIODE(_2833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__A1 (.DIODE(_2833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A1 (.DIODE(_2833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A0 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A1 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__A2 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__B (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A1 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__C (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__A2 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__A1 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__A0 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__B (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A2 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A2 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__B (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__A1 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__A1 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__B (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__A0 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__D (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__D (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__C1 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__C1 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__B (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__B (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__B1 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__B (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__B1 (.DIODE(_2862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__A1 (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__A1 (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__A1 (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__B1 (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__B1 (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__A2 (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__B1 (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__B1 (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__A1 (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__A_N (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__B (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__B (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A1 (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__B (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__B (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__B (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__B (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__B (.DIODE(_2883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__B (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__B1 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A2 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__B2 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__B (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__B1_N (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__A1 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__A1 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__A1 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A1 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__B2 (.DIODE(_2887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__A (.DIODE(_2887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__B2 (.DIODE(_2887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A (.DIODE(_2887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__B2 (.DIODE(_2887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A (.DIODE(_2887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A (.DIODE(_2887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__B2 (.DIODE(_2887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__B2 (.DIODE(_2887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A (.DIODE(_2887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__A (.DIODE(_2888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A (.DIODE(_2888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A (.DIODE(_2888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__A1 (.DIODE(_2888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__A (.DIODE(_2888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__B2 (.DIODE(_2888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__A (.DIODE(_2888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__A1 (.DIODE(_2888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__B2 (.DIODE(_2888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A (.DIODE(_2888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A (.DIODE(_2889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__B1 (.DIODE(_2889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__B (.DIODE(_2889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A1 (.DIODE(_2889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__D (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__A (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__B1 (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__D (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__B (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__D (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__B1 (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A2 (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__D (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__B1 (.DIODE(_2896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__B1 (.DIODE(_2902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A (.DIODE(_2902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__C (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__A (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__A (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__B2 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__B2 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A2 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A2 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__C (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A2 (.DIODE(_2903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__C (.DIODE(_2905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__D (.DIODE(_2905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A (.DIODE(_2905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__C (.DIODE(_2905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__A1 (.DIODE(_2905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A2 (.DIODE(_2905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__B (.DIODE(_2905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__B1 (.DIODE(_2905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__B1 (.DIODE(_2905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__D (.DIODE(_2905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__A (.DIODE(_2916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__A (.DIODE(_2916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A (.DIODE(_2916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A1 (.DIODE(_2916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A (.DIODE(_2916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A1 (.DIODE(_2916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__B2 (.DIODE(_2916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A (.DIODE(_2916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A1 (.DIODE(_2916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__A1 (.DIODE(_2916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__D (.DIODE(_2917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__D (.DIODE(_2917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A (.DIODE(_2917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__A (.DIODE(_2917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__D (.DIODE(_2917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__B2 (.DIODE(_2917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__D (.DIODE(_2917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__B1 (.DIODE(_2917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__B2 (.DIODE(_2917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__B1 (.DIODE(_2917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A (.DIODE(_2921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A (.DIODE(_2921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A (.DIODE(_2921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__A (.DIODE(_2921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__A (.DIODE(_2921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__A (.DIODE(_2921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A (.DIODE(_2921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A (.DIODE(_2921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A (.DIODE(_2921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__A (.DIODE(_2921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__B (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__A (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__A1 (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__A1 (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__A1 (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__B (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__A (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__B2 (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__A (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A1 (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A (.DIODE(_2970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__B (.DIODE(_2970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__A1 (.DIODE(_2984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__A (.DIODE(_2984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A (.DIODE(_2988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__C (.DIODE(_2988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__A (.DIODE(_2988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__C (.DIODE(_2988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__A (.DIODE(_2988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A (.DIODE(_2988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A (.DIODE(_2988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A (.DIODE(_2988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A (.DIODE(_2988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__A1 (.DIODE(_2988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__D (.DIODE(_3001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__D (.DIODE(_3001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__D (.DIODE(_3001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__A2_N (.DIODE(_3001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A2 (.DIODE(_3001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__B1 (.DIODE(_3001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__D (.DIODE(_3001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__B (.DIODE(_3001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__D (.DIODE(_3001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A (.DIODE(_3001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__A0 (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A2_N (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A2_N (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A2_N (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__B (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A1 (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__B (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__A2_N (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__B (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__C (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__B1 (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__B (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__B (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__D (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__A (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__B (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__A (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__A (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__A (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__B1 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__B (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__B (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__B (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A1 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A1 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__B1 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__B1 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__D (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__B1 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A2 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__B (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__B (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__A (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__B2 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__A (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__B2 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__B2 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__A2 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__C (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A2 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__A (.DIODE(_3059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__A (.DIODE(_3059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__B (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__B1_N (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(execute));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(input_val[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(input_val[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(input_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(input_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(input_val[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(input_val[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(input_val[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(input_val[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(reset));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(sel_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(sel_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(sel_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(sel_out[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(sel_out[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A_N (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__A_N (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__A0 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__A0 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__A0 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A0 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout40_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout36_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__B_N (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__D (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__D (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__D_N (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__D (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__D (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__B_N (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__C (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__C (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__D_N (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__C (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__D (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__D_N (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__B_N (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__C (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_output16_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_output17_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_output18_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_output19_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_output20_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_output21_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_output22_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_output23_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_output24_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_output32_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout37_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout39_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__RESET_B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__RESET_B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__RESET_B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__RESET_B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__RESET_B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__RESET_B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__RESET_B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__decap_6 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_841 ();
endmodule

